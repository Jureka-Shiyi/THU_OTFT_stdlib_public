* SPICE NETLIST
***************************************

.SUBCKT INVD2 VSS VDD OUT IN
** N=5 EP=4 IP=0 FDC=12
M0 1 VSS VSS ptft L=4e-05 W=0.0001 $X=-126900 $Y=-172000 $D=0
M1 VDD IN 1 ptft L=1e-05 W=0.0002 $X=-96900 $Y=108000 $D=0
M2 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=-46900 $Y=-172000 $D=0
M3 1 IN VDD ptft L=1e-05 W=0.0002 $X=-46900 $Y=108000 $D=0
M4 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=123100 $Y=-292000 $D=0
M5 VDD IN OUT ptft L=1e-05 W=0.0002 $X=123100 $Y=108000 $D=0
M6 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=173100 $Y=-292000 $D=0
M7 OUT IN VDD ptft L=1e-05 W=0.0002 $X=173100 $Y=108000 $D=0
M8 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=223100 $Y=-292000 $D=0
M9 VDD IN OUT ptft L=1e-05 W=0.0002 $X=223100 $Y=108000 $D=0
M10 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=273100 $Y=-292000 $D=0
M11 OUT IN VDD ptft L=1e-05 W=0.0002 $X=273100 $Y=108000 $D=0
.ENDS
***************************************
