* File: BUFD8.cdl
* Created: Sat Dec 27 13:06:45 2025
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "BUFD8.cdl.pex"
.subckt BUFD8  VSS VDD OUT IN
* 
* IN	IN
* OUT	OUT
* VDD	VDD
* VSS	VSS
XMI5 N_VSS_MI5_d N_VSS_MI5_g N_net3_MI5_s ptft L=4e-05 W=0.0001
XMI5@8 N_VSS_MI5@8_d N_VSS_MI5@8_g N_net3_MI5_s ptft L=4e-05 W=0.0001
XMI5@7 N_VSS_MI5@8_d N_VSS_MI5@7_g N_net3_MI5@7_s ptft L=4e-05 W=0.0001
XMI4 N_net3_MI4_d N_IN_MI4_g N_VDD_MI4_s ptft L=1e-05 W=0.0002
XMI5@6 N_VSS_MI5@6_d N_VSS_MI5@6_g N_net3_MI5@7_s ptft L=4e-05 W=0.0001
XMI4@8 N_net3_MI4@8_d N_IN_MI4@8_g N_VDD_MI4_s ptft L=1e-05 W=0.0002
XMI4@7 N_net3_MI4@8_d N_IN_MI4@7_g N_VDD_MI4@7_s ptft L=1e-05 W=0.0002
XMI5@5 N_VSS_MI5@6_d N_VSS_MI5@5_g N_net3_MI5@5_s ptft L=4e-05 W=0.0001
XMI4@6 N_net3_MI4@6_d N_IN_MI4@6_g N_VDD_MI4@7_s ptft L=1e-05 W=0.0002
XMI5@4 N_VSS_MI5@4_d N_VSS_MI5@4_g N_net3_MI5@5_s ptft L=4e-05 W=0.0001
XMI4@5 N_net3_MI4@6_d N_IN_MI4@5_g N_VDD_MI4@5_s ptft L=1e-05 W=0.0002
XMI4@4 N_net3_MI4@4_d N_IN_MI4@4_g N_VDD_MI4@5_s ptft L=1e-05 W=0.0002
XMI5@3 N_VSS_MI5@4_d N_VSS_MI5@3_g N_net3_MI5@3_s ptft L=4e-05 W=0.0001
XMI4@3 N_net3_MI4@4_d N_IN_MI4@3_g N_VDD_MI4@3_s ptft L=1e-05 W=0.0002
XMI5@2 N_VSS_MI5@2_d N_VSS_MI5@2_g N_net3_MI5@3_s ptft L=4e-05 W=0.0001
XMI4@2 N_net3_MI4@2_d N_IN_MI4@2_g N_VDD_MI4@3_s ptft L=1e-05 W=0.0002
XMI7 N_VSS_MI7_d N_net3_MI7_g N_net1_MI7_s ptft L=1e-05 W=0.0002
XMI6 N_net1_MI6_d N_IN_MI6_g N_VDD_MI6_s ptft L=1e-05 W=0.0002
XMI7@16 N_VSS_MI7_d N_net3_MI7@16_g N_net1_MI7@16_s ptft L=1e-05 W=0.0002
XMI6@16 N_net1_MI6@16_d N_IN_MI6@16_g N_VDD_MI6_s ptft L=1e-05 W=0.0002
XMI7@15 N_VSS_MI7@15_d N_net3_MI7@15_g N_net1_MI7@16_s ptft L=1e-05 W=0.0002
XMI6@15 N_net1_MI6@16_d N_IN_MI6@15_g N_VDD_MI6@15_s ptft L=1e-05 W=0.0002
XMI7@14 N_VSS_MI7@15_d N_net3_MI7@14_g N_net1_MI7@14_s ptft L=1e-05 W=0.0002
XMI6@14 N_net1_MI6@14_d N_IN_MI6@14_g N_VDD_MI6@15_s ptft L=1e-05 W=0.0002
XMI7@13 N_VSS_MI7@13_d N_net3_MI7@13_g N_net1_MI7@14_s ptft L=1e-05 W=0.0002
XMI6@13 N_net1_MI6@14_d N_IN_MI6@13_g N_VDD_MI6@13_s ptft L=1e-05 W=0.0002
XMI7@12 N_VSS_MI7@13_d N_net3_MI7@12_g N_net1_MI7@12_s ptft L=1e-05 W=0.0002
XMI6@12 N_net1_MI6@12_d N_IN_MI6@12_g N_VDD_MI6@13_s ptft L=1e-05 W=0.0002
XMI7@11 N_VSS_MI7@11_d N_net3_MI7@11_g N_net1_MI7@12_s ptft L=1e-05 W=0.0002
XMI6@11 N_net1_MI6@12_d N_IN_MI6@11_g N_VDD_MI6@11_s ptft L=1e-05 W=0.0002
XMI7@10 N_VSS_MI7@11_d N_net3_MI7@10_g N_net1_MI7@10_s ptft L=1e-05 W=0.0002
XMI6@10 N_net1_MI6@10_d N_IN_MI6@10_g N_VDD_MI6@11_s ptft L=1e-05 W=0.0002
XMI7@9 N_VSS_MI7@9_d N_net3_MI7@9_g N_net1_MI7@10_s ptft L=1e-05 W=0.0002
XMI6@9 N_net1_MI6@10_d N_IN_MI6@9_g N_VDD_MI6@9_s ptft L=1e-05 W=0.0002
XMI7@8 N_VSS_MI7@9_d N_net3_MI7@8_g N_net1_MI7@8_s ptft L=1e-05 W=0.0002
XMI6@8 N_net1_MI6@8_d N_IN_MI6@8_g N_VDD_MI6@9_s ptft L=1e-05 W=0.0002
XMI7@7 N_VSS_MI7@7_d N_net3_MI7@7_g N_net1_MI7@8_s ptft L=1e-05 W=0.0002
XMI6@7 N_net1_MI6@8_d N_IN_MI6@7_g N_VDD_MI6@7_s ptft L=1e-05 W=0.0002
XMI7@6 N_VSS_MI7@7_d N_net3_MI7@6_g N_net1_MI7@6_s ptft L=1e-05 W=0.0002
XMI6@6 N_net1_MI6@6_d N_IN_MI6@6_g N_VDD_MI6@7_s ptft L=1e-05 W=0.0002
XMI7@5 N_VSS_MI7@5_d N_net3_MI7@5_g N_net1_MI7@6_s ptft L=1e-05 W=0.0002
XMI6@5 N_net1_MI6@6_d N_IN_MI6@5_g N_VDD_MI6@5_s ptft L=1e-05 W=0.0002
XMI7@4 N_VSS_MI7@5_d N_net3_MI7@4_g N_net1_MI7@4_s ptft L=1e-05 W=0.0002
XMI6@4 N_net1_MI6@4_d N_IN_MI6@4_g N_VDD_MI6@5_s ptft L=1e-05 W=0.0002
XMI7@3 N_VSS_MI7@3_d N_net3_MI7@3_g N_net1_MI7@4_s ptft L=1e-05 W=0.0002
XMI6@3 N_net1_MI6@4_d N_IN_MI6@3_g N_VDD_MI6@3_s ptft L=1e-05 W=0.0002
XMI7@2 N_VSS_MI7@3_d N_net3_MI7@2_g N_net1_MI7@2_s ptft L=1e-05 W=0.0002
XMI6@2 N_net1_MI6@2_d N_IN_MI6@2_g N_VDD_MI6@3_s ptft L=1e-05 W=0.0002
XMI11 N_VSS_MI11_d N_VSS_MI11_g N_net2_MI11_s ptft L=4e-05 W=0.0001
XMI11@8 N_VSS_MI11@8_d N_VSS_MI11@8_g N_net2_MI11_s ptft L=4e-05 W=0.0001
XMI11@7 N_VSS_MI11@8_d N_VSS_MI11@7_g N_net2_MI11@7_s ptft L=4e-05 W=0.0001
XMI9 N_net2_MI9_d N_net1_MI9_g N_VDD_MI9_s ptft L=1e-05 W=0.0002
XMI11@6 N_VSS_MI11@6_d N_VSS_MI11@6_g N_net2_MI11@7_s ptft L=4e-05 W=0.0001
XMI9@8 N_net2_MI9@8_d N_net1_MI9@8_g N_VDD_MI9_s ptft L=1e-05 W=0.0002
XMI9@7 N_net2_MI9@8_d N_net1_MI9@7_g N_VDD_MI9@7_s ptft L=1e-05 W=0.0002
XMI11@5 N_VSS_MI11@6_d N_VSS_MI11@5_g N_net2_MI11@5_s ptft L=4e-05 W=0.0001
XMI9@6 N_net2_MI9@6_d N_net1_MI9@6_g N_VDD_MI9@7_s ptft L=1e-05 W=0.0002
XMI11@4 N_VSS_MI11@4_d N_VSS_MI11@4_g N_net2_MI11@5_s ptft L=4e-05 W=0.0001
XMI9@5 N_net2_MI9@6_d N_net1_MI9@5_g N_VDD_MI9@5_s ptft L=1e-05 W=0.0002
XMI9@4 N_net2_MI9@4_d N_net1_MI9@4_g N_VDD_MI9@5_s ptft L=1e-05 W=0.0002
XMI11@3 N_VSS_MI11@4_d N_VSS_MI11@3_g N_net2_MI11@3_s ptft L=4e-05 W=0.0001
XMI9@3 N_net2_MI9@4_d N_net1_MI9@3_g N_VDD_MI9@3_s ptft L=1e-05 W=0.0002
XMI11@2 N_VSS_MI11@2_d N_VSS_MI11@2_g N_net2_MI11@3_s ptft L=4e-05 W=0.0001
XMI9@2 N_net2_MI9@2_d N_net1_MI9@2_g N_VDD_MI9@3_s ptft L=1e-05 W=0.0002
XMI10 N_VSS_MI10_d N_net2_MI10_g N_OUT_MI10_s ptft L=1e-05 W=0.0002
XMI8 N_OUT_MI8_d N_net1_MI8_g N_VDD_MI8_s ptft L=1e-05 W=0.0002
XMI10@16 N_VSS_MI10_d N_net2_MI10@16_g N_OUT_MI10@16_s ptft L=1e-05 W=0.0002
XMI8@16 N_OUT_MI8@16_d N_net1_MI8@16_g N_VDD_MI8_s ptft L=1e-05 W=0.0002
XMI10@15 N_VSS_MI10@15_d N_net2_MI10@15_g N_OUT_MI10@16_s ptft L=1e-05 W=0.0002
XMI8@15 N_OUT_MI8@16_d N_net1_MI8@15_g N_VDD_MI8@15_s ptft L=1e-05 W=0.0002
XMI10@14 N_VSS_MI10@15_d N_net2_MI10@14_g N_OUT_MI10@14_s ptft L=1e-05 W=0.0002
XMI8@14 N_OUT_MI8@14_d N_net1_MI8@14_g N_VDD_MI8@15_s ptft L=1e-05 W=0.0002
XMI10@13 N_VSS_MI10@13_d N_net2_MI10@13_g N_OUT_MI10@14_s ptft L=1e-05 W=0.0002
XMI8@13 N_OUT_MI8@14_d N_net1_MI8@13_g N_VDD_MI8@13_s ptft L=1e-05 W=0.0002
XMI10@12 N_VSS_MI10@13_d N_net2_MI10@12_g N_OUT_MI10@12_s ptft L=1e-05 W=0.0002
XMI8@12 N_OUT_MI8@12_d N_net1_MI8@12_g N_VDD_MI8@13_s ptft L=1e-05 W=0.0002
XMI10@11 N_VSS_MI10@11_d N_net2_MI10@11_g N_OUT_MI10@12_s ptft L=1e-05 W=0.0002
XMI8@11 N_OUT_MI8@12_d N_net1_MI8@11_g N_VDD_MI8@11_s ptft L=1e-05 W=0.0002
XMI10@10 N_VSS_MI10@11_d N_net2_MI10@10_g N_OUT_MI10@10_s ptft L=1e-05 W=0.0002
XMI8@10 N_OUT_MI8@10_d N_net1_MI8@10_g N_VDD_MI8@11_s ptft L=1e-05 W=0.0002
XMI10@9 N_VSS_MI10@9_d N_net2_MI10@9_g N_OUT_MI10@10_s ptft L=1e-05 W=0.0002
XMI8@9 N_OUT_MI8@10_d N_net1_MI8@9_g N_VDD_MI8@9_s ptft L=1e-05 W=0.0002
XMI10@8 N_VSS_MI10@9_d N_net2_MI10@8_g N_OUT_MI10@8_s ptft L=1e-05 W=0.0002
XMI8@8 N_OUT_MI8@8_d N_net1_MI8@8_g N_VDD_MI8@9_s ptft L=1e-05 W=0.0002
XMI10@7 N_VSS_MI10@7_d N_net2_MI10@7_g N_OUT_MI10@8_s ptft L=1e-05 W=0.0002
XMI8@7 N_OUT_MI8@8_d N_net1_MI8@7_g N_VDD_MI8@7_s ptft L=1e-05 W=0.0002
XMI10@6 N_VSS_MI10@7_d N_net2_MI10@6_g N_OUT_MI10@6_s ptft L=1e-05 W=0.0002
XMI8@6 N_OUT_MI8@6_d N_net1_MI8@6_g N_VDD_MI8@7_s ptft L=1e-05 W=0.0002
XMI10@5 N_VSS_MI10@5_d N_net2_MI10@5_g N_OUT_MI10@6_s ptft L=1e-05 W=0.0002
XMI8@5 N_OUT_MI8@6_d N_net1_MI8@5_g N_VDD_MI8@5_s ptft L=1e-05 W=0.0002
XMI10@4 N_VSS_MI10@5_d N_net2_MI10@4_g N_OUT_MI10@4_s ptft L=1e-05 W=0.0002
XMI8@4 N_OUT_MI8@4_d N_net1_MI8@4_g N_VDD_MI8@5_s ptft L=1e-05 W=0.0002
XMI10@3 N_VSS_MI10@3_d N_net2_MI10@3_g N_OUT_MI10@4_s ptft L=1e-05 W=0.0002
XMI8@3 N_OUT_MI8@4_d N_net1_MI8@3_g N_VDD_MI8@3_s ptft L=1e-05 W=0.0002
XMI10@2 N_VSS_MI10@3_d N_net2_MI10@2_g N_OUT_MI10@2_s ptft L=1e-05 W=0.0002
XMI8@2 N_OUT_MI8@2_d N_net1_MI8@2_g N_VDD_MI8@3_s ptft L=1e-05 W=0.0002
*
.include "BUFD8.cdl.BUFD8.pxi"
*
.ends
*
*
