* SPICE NETLIST
***************************************

.SUBCKT NAND2D1 VSS OUT VDD IN1 IN2
** N=6 EP=5 IP=0 FDC=17
M0 OUT IN1 VDD ptft L=1e-05 W=0.0002 $X=80000 $Y=630000 $D=0
M1 VDD IN1 OUT ptft L=1e-05 W=0.0002 $X=120000 $Y=630000 $D=0
M2 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=140000 $Y=372400 $D=0
M3 OUT IN1 VDD ptft L=1e-05 W=0.0002 $X=160000 $Y=630000 $D=0
M4 VDD IN1 OUT ptft L=1e-05 W=0.0002 $X=200000 $Y=630000 $D=0
M5 1 IN1 VDD ptft L=1e-05 W=0.0002 $X=240000 $Y=630000 $D=0
M6 VDD IN1 1 ptft L=1e-05 W=0.0002 $X=280000 $Y=630000 $D=0
M7 1 IN2 VDD ptft L=1e-05 W=0.0002 $X=320000 $Y=630000 $D=0
M8 VDD IN2 1 ptft L=1e-05 W=0.0002 $X=360000 $Y=630000 $D=0
M9 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=361400 $Y=256600 $D=0
M10 OUT IN2 VDD ptft L=1e-05 W=0.0002 $X=400000 $Y=630000 $D=0
M11 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=401400 $Y=256600 $D=0
M12 VDD IN2 OUT ptft L=1e-05 W=0.0002 $X=440000 $Y=630000 $D=0
M13 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=441400 $Y=256600 $D=0
M14 OUT IN2 VDD ptft L=1e-05 W=0.0002 $X=480000 $Y=630000 $D=0
M15 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=481400 $Y=256600 $D=0
M16 VDD IN2 OUT ptft L=1e-05 W=0.0002 $X=520000 $Y=630000 $D=0
.ENDS
***************************************
