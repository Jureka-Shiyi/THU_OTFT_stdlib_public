* SPICE NETLIST
***************************************

.SUBCKT INVD8 VSS VDD OUT IN
** N=5 EP=4 IP=0 FDC=48
M0 1 VSS VSS ptft L=4e-05 W=0.0001 $X=-606900 $Y=-172000 $D=0
M1 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=-526900 $Y=-172000 $D=0
M2 1 VSS VSS ptft L=4e-05 W=0.0001 $X=-446900 $Y=-172000 $D=0
M3 VDD IN 1 ptft L=1e-05 W=0.0002 $X=-396900 $Y=108000 $D=0
M4 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=-366900 $Y=-172000 $D=0
M5 1 IN VDD ptft L=1e-05 W=0.0002 $X=-346900 $Y=108000 $D=0
M6 VDD IN 1 ptft L=1e-05 W=0.0002 $X=-296900 $Y=108000 $D=0
M7 1 VSS VSS ptft L=4e-05 W=0.0001 $X=-286900 $Y=-172000 $D=0
M8 1 IN VDD ptft L=1e-05 W=0.0002 $X=-246900 $Y=108000 $D=0
M9 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=-206900 $Y=-172000 $D=0
M10 VDD IN 1 ptft L=1e-05 W=0.0002 $X=-196900 $Y=108000 $D=0
M11 1 IN VDD ptft L=1e-05 W=0.0002 $X=-146900 $Y=108000 $D=0
M12 1 VSS VSS ptft L=4e-05 W=0.0001 $X=-126900 $Y=-172000 $D=0
M13 VDD IN 1 ptft L=1e-05 W=0.0002 $X=-96900 $Y=108000 $D=0
M14 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=-46900 $Y=-172000 $D=0
M15 1 IN VDD ptft L=1e-05 W=0.0002 $X=-46900 $Y=108000 $D=0
M16 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=123100 $Y=-292000 $D=0
M17 VDD IN OUT ptft L=1e-05 W=0.0002 $X=123100 $Y=108000 $D=0
M18 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=173100 $Y=-292000 $D=0
M19 OUT IN VDD ptft L=1e-05 W=0.0002 $X=173100 $Y=108000 $D=0
M20 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=223100 $Y=-292000 $D=0
M21 VDD IN OUT ptft L=1e-05 W=0.0002 $X=223100 $Y=108000 $D=0
M22 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=273100 $Y=-292000 $D=0
M23 OUT IN VDD ptft L=1e-05 W=0.0002 $X=273100 $Y=108000 $D=0
M24 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=323100 $Y=-292000 $D=0
M25 VDD IN OUT ptft L=1e-05 W=0.0002 $X=323100 $Y=108000 $D=0
M26 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=373100 $Y=-292000 $D=0
M27 OUT IN VDD ptft L=1e-05 W=0.0002 $X=373100 $Y=108000 $D=0
M28 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=423100 $Y=-292000 $D=0
M29 VDD IN OUT ptft L=1e-05 W=0.0002 $X=423100 $Y=108000 $D=0
M30 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=473100 $Y=-292000 $D=0
M31 OUT IN VDD ptft L=1e-05 W=0.0002 $X=473100 $Y=108000 $D=0
M32 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=523100 $Y=-292000 $D=0
M33 VDD IN OUT ptft L=1e-05 W=0.0002 $X=523100 $Y=108000 $D=0
M34 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=573100 $Y=-292000 $D=0
M35 OUT IN VDD ptft L=1e-05 W=0.0002 $X=573100 $Y=108000 $D=0
M36 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=623100 $Y=-292000 $D=0
M37 VDD IN OUT ptft L=1e-05 W=0.0002 $X=623100 $Y=108000 $D=0
M38 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=673100 $Y=-292000 $D=0
M39 OUT IN VDD ptft L=1e-05 W=0.0002 $X=673100 $Y=108000 $D=0
M40 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=723100 $Y=-292000 $D=0
M41 VDD IN OUT ptft L=1e-05 W=0.0002 $X=723100 $Y=108000 $D=0
M42 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=773100 $Y=-292000 $D=0
M43 OUT IN VDD ptft L=1e-05 W=0.0002 $X=773100 $Y=108000 $D=0
M44 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=823100 $Y=-292000 $D=0
M45 VDD IN OUT ptft L=1e-05 W=0.0002 $X=823100 $Y=108000 $D=0
M46 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=873100 $Y=-292000 $D=0
M47 OUT IN VDD ptft L=1e-05 W=0.0002 $X=873100 $Y=108000 $D=0
.ENDS
***************************************
