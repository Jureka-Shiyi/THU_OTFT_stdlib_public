* SPICE NETLIST
***************************************

.SUBCKT DFFD1 CK D VSS VDD QN Q
** N=26 EP=6 IP=0 FDC=60
M0 VDD 7 4 ptft L=1.8e-05 W=0.00016 $X=540000 $Y=172000 $D=0
M1 VDD CK 5 ptft L=1.8e-05 W=0.00016 $X=540000 $Y=440000 $D=0
M2 VDD D 6 ptft L=1.8e-05 W=0.00016 $X=540000 $Y=708000 $D=0
M3 4 VSS VSS ptft L=1.8e-05 W=4e-05 $X=640000 $Y=70500 $D=0
M4 5 VSS VSS ptft L=1.8e-05 W=4e-05 $X=640000 $Y=338500 $D=0
M5 6 VSS VSS ptft L=1.8e-05 W=4e-05 $X=640000 $Y=606500 $D=0
M6 18 4 VSS ptft L=1.8e-05 W=0.00032 $X=900000 $Y=112000 $D=0
M7 VDD 7 18 ptft L=1.8e-05 W=0.00032 $X=900000 $Y=172000 $D=0
M8 7 5 VSS ptft L=1.8e-05 W=0.00032 $X=900000 $Y=380000 $D=0
M9 VDD CK 7 ptft L=1.8e-05 W=0.00032 $X=900000 $Y=440000 $D=0
M10 10 6 VSS ptft L=1.8e-05 W=0.00032 $X=900000 $Y=648000 $D=0
M11 VDD D 10 ptft L=1.8e-05 W=0.00032 $X=900000 $Y=708000 $D=0
M12 8 7 VDD ptft L=1.8e-05 W=0.00012 $X=1546000 $Y=231000 $D=0
M13 VDD 7 9 ptft L=1.8e-05 W=0.00012 $X=1546000 $Y=615000 $D=0
M14 VSS VSS 8 ptft L=1.8e-05 W=4e-05 $X=1666000 $Y=388500 $D=0
M15 9 VSS VSS ptft L=1.8e-05 W=4e-05 $X=1666000 $Y=457500 $D=0
M16 8 10 VDD ptft L=1.8e-05 W=0.00012 $X=1706000 $Y=231000 $D=0
M17 VDD D 9 ptft L=1.8e-05 W=0.00012 $X=1706000 $Y=615000 $D=0
M18 15 10 VDD ptft L=1.8e-05 W=0.00024 $X=1886000 $Y=231000 $D=0
M19 VDD D 14 ptft L=1.8e-05 W=0.00024 $X=1886000 $Y=615000 $D=0
M20 VSS 8 15 ptft L=1.8e-05 W=0.00048 $X=1926000 $Y=347000 $D=0
M21 14 9 VSS ptft L=1.8e-05 W=0.00048 $X=1926000 $Y=499000 $D=0
M22 15 7 VDD ptft L=1.8e-05 W=0.00024 $X=2166000 $Y=231000 $D=0
M23 VDD 7 14 ptft L=1.8e-05 W=0.00024 $X=2166000 $Y=615000 $D=0
M24 12 17 VDD ptft L=1.8e-05 W=0.00012 $X=2512000 $Y=231000 $D=0
M25 VDD 16 13 ptft L=1.8e-05 W=0.00012 $X=2512000 $Y=615000 $D=0
M26 VSS VSS 12 ptft L=1.8e-05 W=4e-05 $X=2632000 $Y=388500 $D=0
M27 13 VSS VSS ptft L=1.8e-05 W=4e-05 $X=2632000 $Y=457500 $D=0
M28 12 15 VDD ptft L=1.8e-05 W=0.00012 $X=2672000 $Y=231000 $D=0
M29 VDD 14 13 ptft L=1.8e-05 W=0.00012 $X=2672000 $Y=615000 $D=0
M30 16 15 VDD ptft L=1.8e-05 W=0.00024 $X=2852000 $Y=231000 $D=0
M31 VDD 14 17 ptft L=1.8e-05 W=0.00024 $X=2852000 $Y=615000 $D=0
M32 VSS 12 16 ptft L=1.8e-05 W=0.00048 $X=2892000 $Y=347000 $D=0
M33 17 13 VSS ptft L=1.8e-05 W=0.00048 $X=2892000 $Y=499000 $D=0
M34 16 17 VDD ptft L=1.8e-05 W=0.00024 $X=3132000 $Y=231000 $D=0
M35 VDD 16 17 ptft L=1.8e-05 W=0.00024 $X=3132000 $Y=615000 $D=0
M36 19 18 VDD ptft L=1.8e-05 W=0.00012 $X=3646000 $Y=231000 $D=0
M37 VDD 18 20 ptft L=1.8e-05 W=0.00012 $X=3646000 $Y=615000 $D=0
M38 VSS VSS 19 ptft L=1.8e-05 W=4e-05 $X=3766000 $Y=388500 $D=0
M39 20 VSS VSS ptft L=1.8e-05 W=4e-05 $X=3766000 $Y=457500 $D=0
M40 19 16 VDD ptft L=1.8e-05 W=0.00012 $X=3806000 $Y=231000 $D=0
M41 VDD 17 20 ptft L=1.8e-05 W=0.00012 $X=3806000 $Y=615000 $D=0
M42 23 16 VDD ptft L=1.8e-05 W=0.00024 $X=3986000 $Y=231000 $D=0
M43 VDD 17 24 ptft L=1.8e-05 W=0.00024 $X=3986000 $Y=615000 $D=0
M44 VSS 19 23 ptft L=1.8e-05 W=0.00048 $X=4026000 $Y=347000 $D=0
M45 24 20 VSS ptft L=1.8e-05 W=0.00048 $X=4026000 $Y=499000 $D=0
M46 23 18 VDD ptft L=1.8e-05 W=0.00024 $X=4266000 $Y=231000 $D=0
M47 VDD 18 24 ptft L=1.8e-05 W=0.00024 $X=4266000 $Y=615000 $D=0
M48 21 Q VDD ptft L=1.8e-05 W=0.00012 $X=4612000 $Y=231000 $D=0
M49 VDD QN 22 ptft L=1.8e-05 W=0.00012 $X=4612000 $Y=615000 $D=0
M50 VSS VSS 21 ptft L=1.8e-05 W=4e-05 $X=4732000 $Y=388500 $D=0
M51 22 VSS VSS ptft L=1.8e-05 W=4e-05 $X=4732000 $Y=457500 $D=0
M52 21 23 VDD ptft L=1.8e-05 W=0.00012 $X=4772000 $Y=231000 $D=0
M53 VDD 24 22 ptft L=1.8e-05 W=0.00012 $X=4772000 $Y=615000 $D=0
M54 QN 23 VDD ptft L=1.8e-05 W=0.00024 $X=4952000 $Y=231000 $D=0
M55 VDD 24 Q ptft L=1.8e-05 W=0.00024 $X=4952000 $Y=615000 $D=0
M56 VSS 21 QN ptft L=1.8e-05 W=0.00048 $X=4992000 $Y=347000 $D=0
M57 Q 22 VSS ptft L=1.8e-05 W=0.00048 $X=4992000 $Y=499000 $D=0
M58 QN Q VDD ptft L=1.8e-05 W=0.00024 $X=5232000 $Y=231000 $D=0
M59 VDD QN Q ptft L=1.8e-05 W=0.00024 $X=5232000 $Y=615000 $D=0
.ENDS
***************************************
