* SPICE NETLIST
***************************************

.SUBCKT NAND2D2 VSS OUT VDD IN1 IN2
** N=6 EP=5 IP=0 FDC=22
M0 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=10000 $Y=0 $D=0
M1 1 VSS VSS ptft L=1e-05 W=0.0001 $X=30000 $Y=-257600 $D=0
M2 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=50000 $Y=0 $D=0
M3 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=70000 $Y=-257600 $D=0
M4 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=90000 $Y=0 $D=0
M5 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=130000 $Y=0 $D=0
M6 1 IN1 VDD ptft L=1e-05 W=0.0004 $X=170000 $Y=0 $D=0
M7 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=184600 $Y=-386400 $D=0
M8 VDD IN1 1 ptft L=1e-05 W=0.0004 $X=210000 $Y=0 $D=0
M9 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=224600 $Y=-386400 $D=0
M10 1 IN2 VDD ptft L=1e-05 W=0.0004 $X=250000 $Y=0 $D=0
M11 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=264600 $Y=-386400 $D=0
M12 VDD IN2 1 ptft L=1e-05 W=0.0004 $X=290000 $Y=0 $D=0
M13 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=304600 $Y=-386400 $D=0
M14 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=330000 $Y=0 $D=0
M15 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=344600 $Y=-386400 $D=0
M16 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=370000 $Y=0 $D=0
M17 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=384600 $Y=-386400 $D=0
M18 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=410000 $Y=0 $D=0
M19 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=424600 $Y=-386400 $D=0
M20 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=450000 $Y=0 $D=0
M21 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=464600 $Y=-386400 $D=0
.ENDS
***************************************
