* SPICE NETLIST
***************************************

.SUBCKT INVD2 VSS VDD OUT IN
** N=5 EP=4 IP=0 FDC=12
M0 1 VSS VSS ptft L=4e-05 W=0.0001 $X=112000 $Y=300000 $D=0
M1 VDD IN 1 ptft L=1e-05 W=0.0002 $X=142000 $Y=580000 $D=0
M2 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=192000 $Y=300000 $D=0
M3 1 IN VDD ptft L=1e-05 W=0.0002 $X=192000 $Y=580000 $D=0
M4 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=362000 $Y=180000 $D=0
M5 VDD IN OUT ptft L=1e-05 W=0.0002 $X=362000 $Y=580000 $D=0
M6 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=412000 $Y=180000 $D=0
M7 OUT IN VDD ptft L=1e-05 W=0.0002 $X=412000 $Y=580000 $D=0
M8 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=462000 $Y=180000 $D=0
M9 VDD IN OUT ptft L=1e-05 W=0.0002 $X=462000 $Y=580000 $D=0
M10 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=512000 $Y=180000 $D=0
M11 OUT IN VDD ptft L=1e-05 W=0.0002 $X=512000 $Y=580000 $D=0
.ENDS
***************************************
