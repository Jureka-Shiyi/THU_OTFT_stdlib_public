* SPICE NETLIST
***************************************

.SUBCKT NOR2D4 VSS OUT VDD IN2 IN1
** N=8 EP=5 IP=0 FDC=66
M0 2 VSS VSS ptft L=1e-05 W=0.0004 $X=90000 $Y=160000 $D=0
M1 2 IN2 3 ptft L=1e-05 W=0.0002 $X=100000 $Y=310000 $D=0
M2 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=100000 $Y=630000 $D=0
M3 3 IN2 2 ptft L=1e-05 W=0.0002 $X=140000 $Y=310000 $D=0
M4 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=140000 $Y=630000 $D=0
M5 2 IN2 3 ptft L=1e-05 W=0.0002 $X=180000 $Y=310000 $D=0
M6 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=180000 $Y=630000 $D=0
M7 3 IN2 2 ptft L=1e-05 W=0.0002 $X=220000 $Y=310000 $D=0
M8 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=220000 $Y=630000 $D=0
M9 2 IN2 3 ptft L=1e-05 W=0.0002 $X=260000 $Y=310000 $D=0
M10 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=260000 $Y=630000 $D=0
M11 3 IN2 2 ptft L=1e-05 W=0.0002 $X=300000 $Y=310000 $D=0
M12 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=300000 $Y=630000 $D=0
M13 2 IN2 3 ptft L=1e-05 W=0.0002 $X=340000 $Y=310000 $D=0
M14 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=340000 $Y=630000 $D=0
M15 3 IN2 2 ptft L=1e-05 W=0.0002 $X=380000 $Y=310000 $D=0
M16 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=380000 $Y=630000 $D=0
M17 2 IN2 3 ptft L=1e-05 W=0.0002 $X=420000 $Y=310000 $D=0
M18 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=420000 $Y=630000 $D=0
M19 3 IN2 2 ptft L=1e-05 W=0.0002 $X=460000 $Y=310000 $D=0
M20 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=460000 $Y=630000 $D=0
M21 2 IN2 3 ptft L=1e-05 W=0.0002 $X=500000 $Y=310000 $D=0
M22 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=500000 $Y=630000 $D=0
M23 3 IN2 2 ptft L=1e-05 W=0.0002 $X=540000 $Y=310000 $D=0
M24 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=540000 $Y=630000 $D=0
M25 2 IN2 3 ptft L=1e-05 W=0.0002 $X=580000 $Y=310000 $D=0
M26 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=580000 $Y=630000 $D=0
M27 3 IN2 2 ptft L=1e-05 W=0.0002 $X=620000 $Y=310000 $D=0
M28 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=620000 $Y=630000 $D=0
M29 2 IN2 3 ptft L=1e-05 W=0.0002 $X=660000 $Y=310000 $D=0
M30 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=660000 $Y=630000 $D=0
M31 3 IN2 2 ptft L=1e-05 W=0.0002 $X=700000 $Y=310000 $D=0
M32 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=700000 $Y=630000 $D=0
M33 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=810000 $Y=310000 $D=0
M34 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=810000 $Y=630000 $D=0
M35 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=850000 $Y=310000 $D=0
M36 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=850000 $Y=630000 $D=0
M37 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=890000 $Y=310000 $D=0
M38 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=890000 $Y=630000 $D=0
M39 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=930000 $Y=310000 $D=0
M40 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=930000 $Y=630000 $D=0
M41 OUT 2 VSS ptft L=1e-05 W=0.0004 $X=935000 $Y=120000 $D=0
M42 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=970000 $Y=310000 $D=0
M43 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=970000 $Y=630000 $D=0
M44 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=1010000 $Y=310000 $D=0
M45 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=1010000 $Y=630000 $D=0
M46 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=1050000 $Y=310000 $D=0
M47 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=1050000 $Y=630000 $D=0
M48 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=1090000 $Y=310000 $D=0
M49 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=1090000 $Y=630000 $D=0
M50 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=1130000 $Y=310000 $D=0
M51 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=1130000 $Y=630000 $D=0
M52 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=1170000 $Y=310000 $D=0
M53 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=1170000 $Y=630000 $D=0
M54 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=1210000 $Y=310000 $D=0
M55 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=1210000 $Y=630000 $D=0
M56 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=1250000 $Y=310000 $D=0
M57 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=1250000 $Y=630000 $D=0
M58 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=1290000 $Y=310000 $D=0
M59 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=1290000 $Y=630000 $D=0
M60 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=1330000 $Y=310000 $D=0
M61 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=1330000 $Y=630000 $D=0
M62 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=1370000 $Y=310000 $D=0
M63 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=1370000 $Y=630000 $D=0
M64 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=1410000 $Y=310000 $D=0
M65 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=1410000 $Y=630000 $D=0
.ENDS
***************************************
