* SPICE NETLIST
***************************************

.SUBCKT NAND2D2 VSS OUT VDD IN1 IN2
** N=6 EP=5 IP=0 FDC=22
M0 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=80000 $Y=430000 $D=0
M1 1 VSS VSS ptft L=1e-05 W=0.0001 $X=100000 $Y=172400 $D=0
M2 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=120000 $Y=430000 $D=0
M3 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=140000 $Y=172400 $D=0
M4 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=160000 $Y=430000 $D=0
M5 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=200000 $Y=430000 $D=0
M6 1 IN1 VDD ptft L=1e-05 W=0.0004 $X=240000 $Y=430000 $D=0
M7 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=254600 $Y=43600 $D=0
M8 VDD IN1 1 ptft L=1e-05 W=0.0004 $X=280000 $Y=430000 $D=0
M9 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=294600 $Y=43600 $D=0
M10 1 IN2 VDD ptft L=1e-05 W=0.0004 $X=320000 $Y=430000 $D=0
M11 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=334600 $Y=43600 $D=0
M12 VDD IN2 1 ptft L=1e-05 W=0.0004 $X=360000 $Y=430000 $D=0
M13 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=374600 $Y=43600 $D=0
M14 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=400000 $Y=430000 $D=0
M15 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=414600 $Y=43600 $D=0
M16 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=440000 $Y=430000 $D=0
M17 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=454600 $Y=43600 $D=0
M18 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=480000 $Y=430000 $D=0
M19 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=494600 $Y=43600 $D=0
M20 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=520000 $Y=430000 $D=0
M21 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=534600 $Y=43600 $D=0
.ENDS
***************************************
