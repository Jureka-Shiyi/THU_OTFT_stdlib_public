* SPICE NETLIST
***************************************

.SUBCKT NOR2D8 VSS OUT VDD IN2 IN1
** N=8 EP=5 IP=0 FDC=130
M0 2 VSS VSS ptft L=1e-05 W=0.0008 $X=90000 $Y=160000 $D=0
M1 2 IN2 3 ptft L=1e-05 W=0.0002 $X=100000 $Y=310000 $D=0
M2 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=100000 $Y=630000 $D=0
M3 3 IN2 2 ptft L=1e-05 W=0.0002 $X=140000 $Y=310000 $D=0
M4 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=140000 $Y=630000 $D=0
M5 2 IN2 3 ptft L=1e-05 W=0.0002 $X=180000 $Y=310000 $D=0
M6 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=180000 $Y=630000 $D=0
M7 3 IN2 2 ptft L=1e-05 W=0.0002 $X=220000 $Y=310000 $D=0
M8 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=220000 $Y=630000 $D=0
M9 2 IN2 3 ptft L=1e-05 W=0.0002 $X=260000 $Y=310000 $D=0
M10 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=260000 $Y=630000 $D=0
M11 3 IN2 2 ptft L=1e-05 W=0.0002 $X=300000 $Y=310000 $D=0
M12 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=300000 $Y=630000 $D=0
M13 2 IN2 3 ptft L=1e-05 W=0.0002 $X=340000 $Y=310000 $D=0
M14 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=340000 $Y=630000 $D=0
M15 3 IN2 2 ptft L=1e-05 W=0.0002 $X=380000 $Y=310000 $D=0
M16 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=380000 $Y=630000 $D=0
M17 2 IN2 3 ptft L=1e-05 W=0.0002 $X=420000 $Y=310000 $D=0
M18 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=420000 $Y=630000 $D=0
M19 3 IN2 2 ptft L=1e-05 W=0.0002 $X=460000 $Y=310000 $D=0
M20 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=460000 $Y=630000 $D=0
M21 2 IN2 3 ptft L=1e-05 W=0.0002 $X=500000 $Y=310000 $D=0
M22 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=500000 $Y=630000 $D=0
M23 3 IN2 2 ptft L=1e-05 W=0.0002 $X=540000 $Y=310000 $D=0
M24 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=540000 $Y=630000 $D=0
M25 2 IN2 3 ptft L=1e-05 W=0.0002 $X=580000 $Y=310000 $D=0
M26 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=580000 $Y=630000 $D=0
M27 3 IN2 2 ptft L=1e-05 W=0.0002 $X=620000 $Y=310000 $D=0
M28 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=620000 $Y=630000 $D=0
M29 2 IN2 3 ptft L=1e-05 W=0.0002 $X=660000 $Y=310000 $D=0
M30 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=660000 $Y=630000 $D=0
M31 3 IN2 2 ptft L=1e-05 W=0.0002 $X=700000 $Y=310000 $D=0
M32 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=700000 $Y=630000 $D=0
M33 2 IN2 3 ptft L=1e-05 W=0.0002 $X=740000 $Y=310000 $D=0
M34 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=740000 $Y=630000 $D=0
M35 3 IN2 2 ptft L=1e-05 W=0.0002 $X=780000 $Y=310000 $D=0
M36 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=780000 $Y=630000 $D=0
M37 2 IN2 3 ptft L=1e-05 W=0.0002 $X=820000 $Y=310000 $D=0
M38 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=820000 $Y=630000 $D=0
M39 3 IN2 2 ptft L=1e-05 W=0.0002 $X=860000 $Y=310000 $D=0
M40 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=860000 $Y=630000 $D=0
M41 2 IN2 3 ptft L=1e-05 W=0.0002 $X=900000 $Y=310000 $D=0
M42 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=900000 $Y=630000 $D=0
M43 3 IN2 2 ptft L=1e-05 W=0.0002 $X=940000 $Y=310000 $D=0
M44 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=940000 $Y=630000 $D=0
M45 2 IN2 3 ptft L=1e-05 W=0.0002 $X=980000 $Y=310000 $D=0
M46 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=980000 $Y=630000 $D=0
M47 3 IN2 2 ptft L=1e-05 W=0.0002 $X=1020000 $Y=310000 $D=0
M48 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=1020000 $Y=630000 $D=0
M49 2 IN2 3 ptft L=1e-05 W=0.0002 $X=1060000 $Y=310000 $D=0
M50 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=1060000 $Y=630000 $D=0
M51 3 IN2 2 ptft L=1e-05 W=0.0002 $X=1100000 $Y=310000 $D=0
M52 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=1100000 $Y=630000 $D=0
M53 2 IN2 3 ptft L=1e-05 W=0.0002 $X=1140000 $Y=310000 $D=0
M54 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=1140000 $Y=630000 $D=0
M55 3 IN2 2 ptft L=1e-05 W=0.0002 $X=1180000 $Y=310000 $D=0
M56 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=1180000 $Y=630000 $D=0
M57 2 IN2 3 ptft L=1e-05 W=0.0002 $X=1220000 $Y=310000 $D=0
M58 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=1220000 $Y=630000 $D=0
M59 3 IN2 2 ptft L=1e-05 W=0.0002 $X=1260000 $Y=310000 $D=0
M60 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=1260000 $Y=630000 $D=0
M61 2 IN2 3 ptft L=1e-05 W=0.0002 $X=1300000 $Y=310000 $D=0
M62 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=1300000 $Y=630000 $D=0
M63 3 IN2 2 ptft L=1e-05 W=0.0002 $X=1340000 $Y=310000 $D=0
M64 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=1340000 $Y=630000 $D=0
M65 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=1450000 $Y=310000 $D=0
M66 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=1450000 $Y=630000 $D=0
M67 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=1490000 $Y=310000 $D=0
M68 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=1490000 $Y=630000 $D=0
M69 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=1530000 $Y=310000 $D=0
M70 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=1530000 $Y=630000 $D=0
M71 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=1570000 $Y=310000 $D=0
M72 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=1570000 $Y=630000 $D=0
M73 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=1610000 $Y=310000 $D=0
M74 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=1610000 $Y=630000 $D=0
M75 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=1650000 $Y=310000 $D=0
M76 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=1650000 $Y=630000 $D=0
M77 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=1690000 $Y=310000 $D=0
M78 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=1690000 $Y=630000 $D=0
M79 OUT 2 VSS ptft L=1e-05 W=0.0008 $X=1695000 $Y=120000 $D=0
M80 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=1730000 $Y=310000 $D=0
M81 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=1730000 $Y=630000 $D=0
M82 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=1770000 $Y=310000 $D=0
M83 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=1770000 $Y=630000 $D=0
M84 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=1810000 $Y=310000 $D=0
M85 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=1810000 $Y=630000 $D=0
M86 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=1850000 $Y=310000 $D=0
M87 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=1850000 $Y=630000 $D=0
M88 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=1890000 $Y=310000 $D=0
M89 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=1890000 $Y=630000 $D=0
M90 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=1930000 $Y=310000 $D=0
M91 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=1930000 $Y=630000 $D=0
M92 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=1970000 $Y=310000 $D=0
M93 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=1970000 $Y=630000 $D=0
M94 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=2010000 $Y=310000 $D=0
M95 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=2010000 $Y=630000 $D=0
M96 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=2050000 $Y=310000 $D=0
M97 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=2050000 $Y=630000 $D=0
M98 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=2090000 $Y=310000 $D=0
M99 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=2090000 $Y=630000 $D=0
M100 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=2130000 $Y=310000 $D=0
M101 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=2130000 $Y=630000 $D=0
M102 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=2170000 $Y=310000 $D=0
M103 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=2170000 $Y=630000 $D=0
M104 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=2210000 $Y=310000 $D=0
M105 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=2210000 $Y=630000 $D=0
M106 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=2250000 $Y=310000 $D=0
M107 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=2250000 $Y=630000 $D=0
M108 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=2290000 $Y=310000 $D=0
M109 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=2290000 $Y=630000 $D=0
M110 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=2330000 $Y=310000 $D=0
M111 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=2330000 $Y=630000 $D=0
M112 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=2370000 $Y=310000 $D=0
M113 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=2370000 $Y=630000 $D=0
M114 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=2410000 $Y=310000 $D=0
M115 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=2410000 $Y=630000 $D=0
M116 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=2450000 $Y=310000 $D=0
M117 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=2450000 $Y=630000 $D=0
M118 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=2490000 $Y=310000 $D=0
M119 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=2490000 $Y=630000 $D=0
M120 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=2530000 $Y=310000 $D=0
M121 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=2530000 $Y=630000 $D=0
M122 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=2570000 $Y=310000 $D=0
M123 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=2570000 $Y=630000 $D=0
M124 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=2610000 $Y=310000 $D=0
M125 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=2610000 $Y=630000 $D=0
M126 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=2650000 $Y=310000 $D=0
M127 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=2650000 $Y=630000 $D=0
M128 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=2690000 $Y=310000 $D=0
M129 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=2690000 $Y=630000 $D=0
.ENDS
***************************************
