* SPICE NETLIST
***************************************

.SUBCKT NAND2D1 VSS OUT VDD IN1 IN2
** N=6 EP=5 IP=0 FDC=17
M0 OUT IN1 VDD ptft L=1e-05 W=0.0002 $X=10000 $Y=0 $D=0
M1 VDD IN1 OUT ptft L=1e-05 W=0.0002 $X=50000 $Y=0 $D=0
M2 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=70000 $Y=-257600 $D=0
M3 OUT IN1 VDD ptft L=1e-05 W=0.0002 $X=90000 $Y=0 $D=0
M4 VDD IN1 OUT ptft L=1e-05 W=0.0002 $X=130000 $Y=0 $D=0
M5 1 IN1 VDD ptft L=1e-05 W=0.0002 $X=170000 $Y=0 $D=0
M6 VDD IN1 1 ptft L=1e-05 W=0.0002 $X=210000 $Y=0 $D=0
M7 1 IN2 VDD ptft L=1e-05 W=0.0002 $X=250000 $Y=0 $D=0
M8 VDD IN2 1 ptft L=1e-05 W=0.0002 $X=290000 $Y=0 $D=0
M9 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=291400 $Y=-373400 $D=0
M10 OUT IN2 VDD ptft L=1e-05 W=0.0002 $X=330000 $Y=0 $D=0
M11 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=331400 $Y=-373400 $D=0
M12 VDD IN2 OUT ptft L=1e-05 W=0.0002 $X=370000 $Y=0 $D=0
M13 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=371400 $Y=-373400 $D=0
M14 OUT IN2 VDD ptft L=1e-05 W=0.0002 $X=410000 $Y=0 $D=0
M15 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=411400 $Y=-373400 $D=0
M16 VDD IN2 OUT ptft L=1e-05 W=0.0002 $X=450000 $Y=0 $D=0
.ENDS
***************************************
