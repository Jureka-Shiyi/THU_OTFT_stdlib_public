* SPICE NETLIST
***************************************

.SUBCKT INVD8 VSS VDD OUT IN
** N=5 EP=4 IP=0 FDC=48
M0 1 VSS VSS ptft L=4e-05 W=0.0001 $X=80000 $Y=300000 $D=0
M1 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=160000 $Y=300000 $D=0
M2 1 VSS VSS ptft L=4e-05 W=0.0001 $X=240000 $Y=300000 $D=0
M3 VDD IN 1 ptft L=1e-05 W=0.0002 $X=290000 $Y=580000 $D=0
M4 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=320000 $Y=300000 $D=0
M5 1 IN VDD ptft L=1e-05 W=0.0002 $X=340000 $Y=580000 $D=0
M6 VDD IN 1 ptft L=1e-05 W=0.0002 $X=390000 $Y=580000 $D=0
M7 1 VSS VSS ptft L=4e-05 W=0.0001 $X=400000 $Y=300000 $D=0
M8 1 IN VDD ptft L=1e-05 W=0.0002 $X=440000 $Y=580000 $D=0
M9 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=480000 $Y=300000 $D=0
M10 VDD IN 1 ptft L=1e-05 W=0.0002 $X=490000 $Y=580000 $D=0
M11 1 IN VDD ptft L=1e-05 W=0.0002 $X=540000 $Y=580000 $D=0
M12 1 VSS VSS ptft L=4e-05 W=0.0001 $X=560000 $Y=300000 $D=0
M13 VDD IN 1 ptft L=1e-05 W=0.0002 $X=590000 $Y=580000 $D=0
M14 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=640000 $Y=300000 $D=0
M15 1 IN VDD ptft L=1e-05 W=0.0002 $X=640000 $Y=580000 $D=0
M16 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=810000 $Y=180000 $D=0
M17 VDD IN OUT ptft L=1e-05 W=0.0002 $X=810000 $Y=580000 $D=0
M18 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=860000 $Y=180000 $D=0
M19 OUT IN VDD ptft L=1e-05 W=0.0002 $X=860000 $Y=580000 $D=0
M20 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=910000 $Y=180000 $D=0
M21 VDD IN OUT ptft L=1e-05 W=0.0002 $X=910000 $Y=580000 $D=0
M22 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=960000 $Y=180000 $D=0
M23 OUT IN VDD ptft L=1e-05 W=0.0002 $X=960000 $Y=580000 $D=0
M24 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1010000 $Y=180000 $D=0
M25 VDD IN OUT ptft L=1e-05 W=0.0002 $X=1010000 $Y=580000 $D=0
M26 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1060000 $Y=180000 $D=0
M27 OUT IN VDD ptft L=1e-05 W=0.0002 $X=1060000 $Y=580000 $D=0
M28 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1110000 $Y=180000 $D=0
M29 VDD IN OUT ptft L=1e-05 W=0.0002 $X=1110000 $Y=580000 $D=0
M30 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1160000 $Y=180000 $D=0
M31 OUT IN VDD ptft L=1e-05 W=0.0002 $X=1160000 $Y=580000 $D=0
M32 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1210000 $Y=180000 $D=0
M33 VDD IN OUT ptft L=1e-05 W=0.0002 $X=1210000 $Y=580000 $D=0
M34 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1260000 $Y=180000 $D=0
M35 OUT IN VDD ptft L=1e-05 W=0.0002 $X=1260000 $Y=580000 $D=0
M36 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1310000 $Y=180000 $D=0
M37 VDD IN OUT ptft L=1e-05 W=0.0002 $X=1310000 $Y=580000 $D=0
M38 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1360000 $Y=180000 $D=0
M39 OUT IN VDD ptft L=1e-05 W=0.0002 $X=1360000 $Y=580000 $D=0
M40 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1410000 $Y=180000 $D=0
M41 VDD IN OUT ptft L=1e-05 W=0.0002 $X=1410000 $Y=580000 $D=0
M42 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1460000 $Y=180000 $D=0
M43 OUT IN VDD ptft L=1e-05 W=0.0002 $X=1460000 $Y=580000 $D=0
M44 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1510000 $Y=180000 $D=0
M45 VDD IN OUT ptft L=1e-05 W=0.0002 $X=1510000 $Y=580000 $D=0
M46 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1560000 $Y=180000 $D=0
M47 OUT IN VDD ptft L=1e-05 W=0.0002 $X=1560000 $Y=580000 $D=0
.ENDS
***************************************
