* File: OR2D1.cdl
* Created: Wed Jan 15 19:04:35 2025
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "/data/zhengyj/OTFT_stdlib/subckts/OR2D1.cdl.pex"
.subckt OR2D1  IN1 IN2 VSS VDD OUT
* 
* OUT	OUT
* VDD	VDD
* VSS	VSS
* IN2	IN2
* IN1	IN1
XMI5 N_OUT_MI5_d N_net12_MI5_g N_VSS_MI5_s ntft L=4e-06 W=4e-05
XMI3 N_net12_MI3_d N_IN1_MI3_g N_VSS_MI3_s ntft L=4e-06 W=2e-05
XMI4 N_net12_MI4_d N_IN2_MI4_g N_VSS_MI4_s ntft L=4e-06 W=2e-05
XMI6 N_net12_MI6_d N_IN2_MI6_g net11 ptft L=4e-06 W=2e-05
XMI0 net11 N_IN1_MI0_g N_VDD_MI0_s ptft L=4e-06 W=2e-05
XMI7 N_OUT_MI7_d N_net12_MI7_g N_VDD_MI7_s ptft L=4e-06 W=2e-05
c_129 net11 0 0.143191f
*
.include "/data/zhengyj/OTFT_stdlib/subckts/OR2D1.cdl.OR2D1.pxi"
*
.ends
*
*
