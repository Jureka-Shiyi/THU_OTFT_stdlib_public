
*************************************************************
*** EsimFPD Model ver: 2021.10.hf1                        ***
***       Built at: 12/30/2021 20:15                      ***
***   (C) Copyright 2021 Huada Empyrean Software Co.      ***
*************************************************************
.model otft_ito_2  pmos
+ level= 62             
+ version= 1              
+ capmod= 0              
+ shmod= 0              
+ isubmod= 0              
+ idsmod= 1              
+ vtmod= 1              
+ diblmod= 1              
+ acm= 0              
+ wmin= 0.0015         
+ wmax= 0.0015         
+ lmin= 5e-05          
+ lmax= 5e-05          
+ zeroc= 0              
+ cornermod= 0              
+ binmod= 0              
+ tox= 1e-07          
+ eps= 11.7           
+ epsi= 2.82           
+ ld= 0              
+ wd= 0              
+ ldif= 0              
+ hdif= 0              
+ wmlt= 1              
+ lmlt= 1              
+ xw= 0              
+ xl= 0              
+ xj= 1.5e-07        
+ del= 0              
+ vto= -0.266616      
+ von= 0              
+ vfb= 0.310911       
+ vsi= 2.0402         
+ vst= 1.65234        
+ at= 2.40489e-08    
+ bt= 1.55402e-06    
+ dvt= 0.1            
+ cgso= 0              
+ cgdo= 0              
+ etac0= 7              
+ etac00= 0              
+ mc= 3              
+ kss= 0              
+ rsx= 0              
+ rdx= 0              
+ eta= 2.78239        
+ delta= 1.61408        
+ mus= 0.0450607      
+ mu0= 81.7907        
+ mu1= 0.00112029     
+ mmu= 1.13725        
+ meta= 1              
+ theta= 1e-09          
+ ad= 593588         
+ ag= 1.1448e+07     
+ dd= 1.68467e-06    
+ dg= 8.73514e-08    
+ blk= 7.47963e-05    
+ i0= 0.811998       
+ eb= 0.880774       
+ i00= 150            
+ alphasat= 0.929645       
+ lasat= 2.5e-07        
+ me= 2.5            
+ mss= 3              
+ vmax= 40000          
+ lambda= 0.048          
+ ls= 3.5e-08        
+ vp= 0.2            
+ lkink= 5e-05          
+ mk= 1              
+ vkink= 33.4701        
+ tnom= 27             
+ dvto= 0              
+ dmu1= 0              
+ dasat= 0              
+ kt1= 0              
+ teta= 0              
+ ute= 0              
+ mus1= 0              
+ vat= 0              
+ kat= 0              
+ kbt= 0              
+ prt= 0              
+ kasat= 0              
+ ki0= 0              
+ ki00= 0              
+ rth0= 0              
+ cth0= 0              
+ intdsnod= 0              
+ rsh= 0              
+ rd= 0              
+ rs= 0              
+ rdc= 0              
+ rsc= 0              




************************************************************
****                                     Data        Model
**** Eff. Mobility(cm2/volt/sec)      0.31777     0.723362
****                      Vth(V)     -1.41457     -1.40463
****  Sub-Threshold Slope(V/dec)     0.447397     0.456119
****          Ion(A) @ Vgs = 10V  1.38455e-05  2.12945e-05
****        Ioff(A) @ Vgs = -10V    6.562e-12  2.23731e-12
************************************************************

