* File: NOR2D1.cdl
* Created: Sat Aug 17 14:54:54 2024
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "/data/zhengyj/OTFT_stdlib/subckts/NOR2D1.cdl.pex"
.subckt NOR2D1  IN1 IN2 VSS VDD OUT
* 
* OUT	OUT
* VDD	VDD
* VSS	VSS
* IN2	IN2
* IN1	IN1
XMI0 N_OUT_MI0_d N_IN1_MI0_g N_VSS_MI0_s ntft L=4e-06 W=2e-05
XMI1 N_OUT_MI1_d N_IN2_MI1_g N_VSS_MI1_s ntft L=4e-06 W=2e-05
XMI7 N_OUT_MI7_d N_IN2_MI7_g net1 ptft L=4e-06 W=2e-05
XMI6 net1 N_IN1_MI6_g N_VDD_MI6_s ptft L=4e-06 W=2e-05
c_73 net1 0 0.245868f
*
.include "/data/zhengyj/OTFT_stdlib/subckts/NOR2D1.cdl.NOR2D1.pxi"
*
.ends
*
*
