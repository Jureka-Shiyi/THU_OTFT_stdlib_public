* SPICE NETLIST
***************************************

.SUBCKT BUFD8 VSS VDD OUT IN
** N=7 EP=4 IP=0 FDC=96
M0 1 VSS VSS ptft L=4e-05 W=0.0001 $X=80000 $Y=300000 $D=0
M1 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=160000 $Y=300000 $D=0
M2 1 VSS VSS ptft L=4e-05 W=0.0001 $X=240000 $Y=300000 $D=0
M3 VDD IN 1 ptft L=1e-05 W=0.0002 $X=290000 $Y=580000 $D=0
M4 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=320000 $Y=300000 $D=0
M5 1 IN VDD ptft L=1e-05 W=0.0002 $X=340000 $Y=580000 $D=0
M6 VDD IN 1 ptft L=1e-05 W=0.0002 $X=390000 $Y=580000 $D=0
M7 1 VSS VSS ptft L=4e-05 W=0.0001 $X=400000 $Y=300000 $D=0
M8 1 IN VDD ptft L=1e-05 W=0.0002 $X=440000 $Y=580000 $D=0
M9 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=480000 $Y=300000 $D=0
M10 VDD IN 1 ptft L=1e-05 W=0.0002 $X=490000 $Y=580000 $D=0
M11 1 IN VDD ptft L=1e-05 W=0.0002 $X=540000 $Y=580000 $D=0
M12 1 VSS VSS ptft L=4e-05 W=0.0001 $X=560000 $Y=300000 $D=0
M13 VDD IN 1 ptft L=1e-05 W=0.0002 $X=590000 $Y=580000 $D=0
M14 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=640000 $Y=300000 $D=0
M15 1 IN VDD ptft L=1e-05 W=0.0002 $X=640000 $Y=580000 $D=0
M16 VSS 1 3 ptft L=1e-05 W=0.0002 $X=810000 $Y=180000 $D=0
M17 VDD IN 3 ptft L=1e-05 W=0.0002 $X=810000 $Y=580000 $D=0
M18 3 1 VSS ptft L=1e-05 W=0.0002 $X=860000 $Y=180000 $D=0
M19 3 IN VDD ptft L=1e-05 W=0.0002 $X=860000 $Y=580000 $D=0
M20 VSS 1 3 ptft L=1e-05 W=0.0002 $X=910000 $Y=180000 $D=0
M21 VDD IN 3 ptft L=1e-05 W=0.0002 $X=910000 $Y=580000 $D=0
M22 3 1 VSS ptft L=1e-05 W=0.0002 $X=960000 $Y=180000 $D=0
M23 3 IN VDD ptft L=1e-05 W=0.0002 $X=960000 $Y=580000 $D=0
M24 VSS 1 3 ptft L=1e-05 W=0.0002 $X=1010000 $Y=180000 $D=0
M25 VDD IN 3 ptft L=1e-05 W=0.0002 $X=1010000 $Y=580000 $D=0
M26 3 1 VSS ptft L=1e-05 W=0.0002 $X=1060000 $Y=180000 $D=0
M27 3 IN VDD ptft L=1e-05 W=0.0002 $X=1060000 $Y=580000 $D=0
M28 VSS 1 3 ptft L=1e-05 W=0.0002 $X=1110000 $Y=180000 $D=0
M29 VDD IN 3 ptft L=1e-05 W=0.0002 $X=1110000 $Y=580000 $D=0
M30 3 1 VSS ptft L=1e-05 W=0.0002 $X=1160000 $Y=180000 $D=0
M31 3 IN VDD ptft L=1e-05 W=0.0002 $X=1160000 $Y=580000 $D=0
M32 VSS 1 3 ptft L=1e-05 W=0.0002 $X=1210000 $Y=180000 $D=0
M33 VDD IN 3 ptft L=1e-05 W=0.0002 $X=1210000 $Y=580000 $D=0
M34 3 1 VSS ptft L=1e-05 W=0.0002 $X=1260000 $Y=180000 $D=0
M35 3 IN VDD ptft L=1e-05 W=0.0002 $X=1260000 $Y=580000 $D=0
M36 VSS 1 3 ptft L=1e-05 W=0.0002 $X=1310000 $Y=180000 $D=0
M37 VDD IN 3 ptft L=1e-05 W=0.0002 $X=1310000 $Y=580000 $D=0
M38 3 1 VSS ptft L=1e-05 W=0.0002 $X=1360000 $Y=180000 $D=0
M39 3 IN VDD ptft L=1e-05 W=0.0002 $X=1360000 $Y=580000 $D=0
M40 VSS 1 3 ptft L=1e-05 W=0.0002 $X=1410000 $Y=180000 $D=0
M41 VDD IN 3 ptft L=1e-05 W=0.0002 $X=1410000 $Y=580000 $D=0
M42 3 1 VSS ptft L=1e-05 W=0.0002 $X=1460000 $Y=180000 $D=0
M43 3 IN VDD ptft L=1e-05 W=0.0002 $X=1460000 $Y=580000 $D=0
M44 VSS 1 3 ptft L=1e-05 W=0.0002 $X=1510000 $Y=180000 $D=0
M45 VDD IN 3 ptft L=1e-05 W=0.0002 $X=1510000 $Y=580000 $D=0
M46 3 1 VSS ptft L=1e-05 W=0.0002 $X=1560000 $Y=180000 $D=0
M47 3 IN VDD ptft L=1e-05 W=0.0002 $X=1560000 $Y=580000 $D=0
M48 4 VSS VSS ptft L=4e-05 W=0.0001 $X=1720000 $Y=300000 $D=0
M49 VSS VSS 4 ptft L=4e-05 W=0.0001 $X=1800000 $Y=300000 $D=0
M50 4 VSS VSS ptft L=4e-05 W=0.0001 $X=1880000 $Y=300000 $D=0
M51 VDD 3 4 ptft L=1e-05 W=0.0002 $X=1930000 $Y=580000 $D=0
M52 VSS VSS 4 ptft L=4e-05 W=0.0001 $X=1960000 $Y=300000 $D=0
M53 4 3 VDD ptft L=1e-05 W=0.0002 $X=1980000 $Y=580000 $D=0
M54 VDD 3 4 ptft L=1e-05 W=0.0002 $X=2030000 $Y=580000 $D=0
M55 4 VSS VSS ptft L=4e-05 W=0.0001 $X=2040000 $Y=300000 $D=0
M56 4 3 VDD ptft L=1e-05 W=0.0002 $X=2080000 $Y=580000 $D=0
M57 VSS VSS 4 ptft L=4e-05 W=0.0001 $X=2120000 $Y=300000 $D=0
M58 VDD 3 4 ptft L=1e-05 W=0.0002 $X=2130000 $Y=580000 $D=0
M59 4 3 VDD ptft L=1e-05 W=0.0002 $X=2180000 $Y=580000 $D=0
M60 4 VSS VSS ptft L=4e-05 W=0.0001 $X=2200000 $Y=300000 $D=0
M61 VDD 3 4 ptft L=1e-05 W=0.0002 $X=2230000 $Y=580000 $D=0
M62 VSS VSS 4 ptft L=4e-05 W=0.0001 $X=2280000 $Y=300000 $D=0
M63 4 3 VDD ptft L=1e-05 W=0.0002 $X=2280000 $Y=580000 $D=0
M64 VSS 4 OUT ptft L=1e-05 W=0.0002 $X=2450000 $Y=180000 $D=0
M65 VDD 3 OUT ptft L=1e-05 W=0.0002 $X=2450000 $Y=580000 $D=0
M66 OUT 4 VSS ptft L=1e-05 W=0.0002 $X=2500000 $Y=180000 $D=0
M67 OUT 3 VDD ptft L=1e-05 W=0.0002 $X=2500000 $Y=580000 $D=0
M68 VSS 4 OUT ptft L=1e-05 W=0.0002 $X=2550000 $Y=180000 $D=0
M69 VDD 3 OUT ptft L=1e-05 W=0.0002 $X=2550000 $Y=580000 $D=0
M70 OUT 4 VSS ptft L=1e-05 W=0.0002 $X=2600000 $Y=180000 $D=0
M71 OUT 3 VDD ptft L=1e-05 W=0.0002 $X=2600000 $Y=580000 $D=0
M72 VSS 4 OUT ptft L=1e-05 W=0.0002 $X=2650000 $Y=180000 $D=0
M73 VDD 3 OUT ptft L=1e-05 W=0.0002 $X=2650000 $Y=580000 $D=0
M74 OUT 4 VSS ptft L=1e-05 W=0.0002 $X=2700000 $Y=180000 $D=0
M75 OUT 3 VDD ptft L=1e-05 W=0.0002 $X=2700000 $Y=580000 $D=0
M76 VSS 4 OUT ptft L=1e-05 W=0.0002 $X=2750000 $Y=180000 $D=0
M77 VDD 3 OUT ptft L=1e-05 W=0.0002 $X=2750000 $Y=580000 $D=0
M78 OUT 4 VSS ptft L=1e-05 W=0.0002 $X=2800000 $Y=180000 $D=0
M79 OUT 3 VDD ptft L=1e-05 W=0.0002 $X=2800000 $Y=580000 $D=0
M80 VSS 4 OUT ptft L=1e-05 W=0.0002 $X=2850000 $Y=180000 $D=0
M81 VDD 3 OUT ptft L=1e-05 W=0.0002 $X=2850000 $Y=580000 $D=0
M82 OUT 4 VSS ptft L=1e-05 W=0.0002 $X=2900000 $Y=180000 $D=0
M83 OUT 3 VDD ptft L=1e-05 W=0.0002 $X=2900000 $Y=580000 $D=0
M84 VSS 4 OUT ptft L=1e-05 W=0.0002 $X=2950000 $Y=180000 $D=0
M85 VDD 3 OUT ptft L=1e-05 W=0.0002 $X=2950000 $Y=580000 $D=0
M86 OUT 4 VSS ptft L=1e-05 W=0.0002 $X=3000000 $Y=180000 $D=0
M87 OUT 3 VDD ptft L=1e-05 W=0.0002 $X=3000000 $Y=580000 $D=0
M88 VSS 4 OUT ptft L=1e-05 W=0.0002 $X=3050000 $Y=180000 $D=0
M89 VDD 3 OUT ptft L=1e-05 W=0.0002 $X=3050000 $Y=580000 $D=0
M90 OUT 4 VSS ptft L=1e-05 W=0.0002 $X=3100000 $Y=180000 $D=0
M91 OUT 3 VDD ptft L=1e-05 W=0.0002 $X=3100000 $Y=580000 $D=0
M92 VSS 4 OUT ptft L=1e-05 W=0.0002 $X=3150000 $Y=180000 $D=0
M93 VDD 3 OUT ptft L=1e-05 W=0.0002 $X=3150000 $Y=580000 $D=0
M94 OUT 4 VSS ptft L=1e-05 W=0.0002 $X=3200000 $Y=180000 $D=0
M95 OUT 3 VDD ptft L=1e-05 W=0.0002 $X=3200000 $Y=580000 $D=0
.ENDS
***************************************
