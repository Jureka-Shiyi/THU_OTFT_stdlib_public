* File: INVD8.cdl
* Created: Mon Dec 22 20:56:18 2025
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "/data/zhengyj/OTFT_stdlib/subckts_cdl/INVD8.cdl.pex"
.subckt INVD8  VSS VDD OUT IN
* 
* IN	IN
* OUT	OUT
* VDD	VDD
* VSS	VSS
XMI5 N_VSS_MI5_d N_VSS_MI5_g N_net10_MI5_s ptft L=4e-05 W=0.0001
XMI5@8 N_VSS_MI5@8_d N_VSS_MI5@8_g N_net10_MI5_s ptft L=4e-05 W=0.0001
XMI5@7 N_VSS_MI5@8_d N_VSS_MI5@7_g N_net10_MI5@7_s ptft L=4e-05 W=0.0001
XMI4 N_net10_MI4_d N_IN_MI4_g N_VDD_MI4_s ptft L=1e-05 W=0.0002
XMI5@6 N_VSS_MI5@6_d N_VSS_MI5@6_g N_net10_MI5@7_s ptft L=4e-05 W=0.0001
XMI4@8 N_net10_MI4@8_d N_IN_MI4@8_g N_VDD_MI4_s ptft L=1e-05 W=0.0002
XMI4@7 N_net10_MI4@8_d N_IN_MI4@7_g N_VDD_MI4@7_s ptft L=1e-05 W=0.0002
XMI5@5 N_VSS_MI5@6_d N_VSS_MI5@5_g N_net10_MI5@5_s ptft L=4e-05 W=0.0001
XMI4@6 N_net10_MI4@6_d N_IN_MI4@6_g N_VDD_MI4@7_s ptft L=1e-05 W=0.0002
XMI5@4 N_VSS_MI5@4_d N_VSS_MI5@4_g N_net10_MI5@5_s ptft L=4e-05 W=0.0001
XMI4@5 N_net10_MI4@6_d N_IN_MI4@5_g N_VDD_MI4@5_s ptft L=1e-05 W=0.0002
XMI4@4 N_net10_MI4@4_d N_IN_MI4@4_g N_VDD_MI4@5_s ptft L=1e-05 W=0.0002
XMI5@3 N_VSS_MI5@4_d N_VSS_MI5@3_g N_net10_MI5@3_s ptft L=4e-05 W=0.0001
XMI4@3 N_net10_MI4@4_d N_IN_MI4@3_g N_VDD_MI4@3_s ptft L=1e-05 W=0.0002
XMI5@2 N_VSS_MI5@2_d N_VSS_MI5@2_g N_net10_MI5@3_s ptft L=4e-05 W=0.0001
XMI4@2 N_net10_MI4@2_d N_IN_MI4@2_g N_VDD_MI4@3_s ptft L=1e-05 W=0.0002
XMI7 N_VSS_MI7_d N_net10_MI7_g N_OUT_MI7_s ptft L=1e-05 W=0.0002
XMI6 N_OUT_MI6_d N_IN_MI6_g N_VDD_MI6_s ptft L=1e-05 W=0.0002
XMI7@16 N_VSS_MI7_d N_net10_MI7@16_g N_OUT_MI7@16_s ptft L=1e-05 W=0.0002
XMI6@16 N_OUT_MI6@16_d N_IN_MI6@16_g N_VDD_MI6_s ptft L=1e-05 W=0.0002
XMI7@15 N_VSS_MI7@15_d N_net10_MI7@15_g N_OUT_MI7@16_s ptft L=1e-05 W=0.0002
XMI6@15 N_OUT_MI6@16_d N_IN_MI6@15_g N_VDD_MI6@15_s ptft L=1e-05 W=0.0002
XMI7@14 N_VSS_MI7@15_d N_net10_MI7@14_g N_OUT_MI7@14_s ptft L=1e-05 W=0.0002
XMI6@14 N_OUT_MI6@14_d N_IN_MI6@14_g N_VDD_MI6@15_s ptft L=1e-05 W=0.0002
XMI7@13 N_VSS_MI7@13_d N_net10_MI7@13_g N_OUT_MI7@14_s ptft L=1e-05 W=0.0002
XMI6@13 N_OUT_MI6@14_d N_IN_MI6@13_g N_VDD_MI6@13_s ptft L=1e-05 W=0.0002
XMI7@12 N_VSS_MI7@13_d N_net10_MI7@12_g N_OUT_MI7@12_s ptft L=1e-05 W=0.0002
XMI6@12 N_OUT_MI6@12_d N_IN_MI6@12_g N_VDD_MI6@13_s ptft L=1e-05 W=0.0002
XMI7@11 N_VSS_MI7@11_d N_net10_MI7@11_g N_OUT_MI7@12_s ptft L=1e-05 W=0.0002
XMI6@11 N_OUT_MI6@12_d N_IN_MI6@11_g N_VDD_MI6@11_s ptft L=1e-05 W=0.0002
XMI7@10 N_VSS_MI7@11_d N_net10_MI7@10_g N_OUT_MI7@10_s ptft L=1e-05 W=0.0002
XMI6@10 N_OUT_MI6@10_d N_IN_MI6@10_g N_VDD_MI6@11_s ptft L=1e-05 W=0.0002
XMI7@9 N_VSS_MI7@9_d N_net10_MI7@9_g N_OUT_MI7@10_s ptft L=1e-05 W=0.0002
XMI6@9 N_OUT_MI6@10_d N_IN_MI6@9_g N_VDD_MI6@9_s ptft L=1e-05 W=0.0002
XMI7@8 N_VSS_MI7@9_d N_net10_MI7@8_g N_OUT_MI7@8_s ptft L=1e-05 W=0.0002
XMI6@8 N_OUT_MI6@8_d N_IN_MI6@8_g N_VDD_MI6@9_s ptft L=1e-05 W=0.0002
XMI7@7 N_VSS_MI7@7_d N_net10_MI7@7_g N_OUT_MI7@8_s ptft L=1e-05 W=0.0002
XMI6@7 N_OUT_MI6@8_d N_IN_MI6@7_g N_VDD_MI6@7_s ptft L=1e-05 W=0.0002
XMI7@6 N_VSS_MI7@7_d N_net10_MI7@6_g N_OUT_MI7@6_s ptft L=1e-05 W=0.0002
XMI6@6 N_OUT_MI6@6_d N_IN_MI6@6_g N_VDD_MI6@7_s ptft L=1e-05 W=0.0002
XMI7@5 N_VSS_MI7@5_d N_net10_MI7@5_g N_OUT_MI7@6_s ptft L=1e-05 W=0.0002
XMI6@5 N_OUT_MI6@6_d N_IN_MI6@5_g N_VDD_MI6@5_s ptft L=1e-05 W=0.0002
XMI7@4 N_VSS_MI7@5_d N_net10_MI7@4_g N_OUT_MI7@4_s ptft L=1e-05 W=0.0002
XMI6@4 N_OUT_MI6@4_d N_IN_MI6@4_g N_VDD_MI6@5_s ptft L=1e-05 W=0.0002
XMI7@3 N_VSS_MI7@3_d N_net10_MI7@3_g N_OUT_MI7@4_s ptft L=1e-05 W=0.0002
XMI6@3 N_OUT_MI6@4_d N_IN_MI6@3_g N_VDD_MI6@3_s ptft L=1e-05 W=0.0002
XMI7@2 N_VSS_MI7@3_d N_net10_MI7@2_g N_OUT_MI7@2_s ptft L=1e-05 W=0.0002
XMI6@2 N_OUT_MI6@2_d N_IN_MI6@2_g N_VDD_MI6@3_s ptft L=1e-05 W=0.0002
*
.include "/data/zhengyj/OTFT_stdlib/subckts_cdl/INVD8.cdl.INVD8.pxi"
*
.ends
*
*
