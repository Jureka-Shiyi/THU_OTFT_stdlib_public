* SPICE NETLIST
***************************************

.SUBCKT NAND2D8 VSS OUT VDD IN1 IN2
** N=6 EP=5 IP=0 FDC=88
M0 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=-710000 $Y=0 $D=0
M1 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=-670000 $Y=0 $D=0
M2 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=-630000 $Y=0 $D=0
M3 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=-590000 $Y=0 $D=0
M4 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=-550000 $Y=0 $D=0
M5 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=-510000 $Y=0 $D=0
M6 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=-470000 $Y=0 $D=0
M7 1 VSS VSS ptft L=1e-05 W=0.0001 $X=-464600 $Y=-257600 $D=0
M8 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=-430000 $Y=0 $D=0
M9 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=-424600 $Y=-257600 $D=0
M10 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=-390000 $Y=0 $D=0
M11 1 VSS VSS ptft L=1e-05 W=0.0001 $X=-384600 $Y=-257600 $D=0
M12 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=-350000 $Y=0 $D=0
M13 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=-344600 $Y=-257600 $D=0
M14 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=-310000 $Y=0 $D=0
M15 1 VSS VSS ptft L=1e-05 W=0.0001 $X=-304600 $Y=-257600 $D=0
M16 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=-270000 $Y=0 $D=0
M17 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=-264600 $Y=-257600 $D=0
M18 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=-230000 $Y=0 $D=0
M19 1 VSS VSS ptft L=1e-05 W=0.0001 $X=-224600 $Y=-257600 $D=0
M20 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=-190000 $Y=0 $D=0
M21 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=-184600 $Y=-257600 $D=0
M22 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=-150000 $Y=0 $D=0
M23 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=-110000 $Y=0 $D=0
M24 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=-70000 $Y=-386400 $D=0
M25 1 IN1 VDD ptft L=1e-05 W=0.0004 $X=-70000 $Y=0 $D=0
M26 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=-30000 $Y=-386400 $D=0
M27 VDD IN1 1 ptft L=1e-05 W=0.0004 $X=-30000 $Y=0 $D=0
M28 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=10000 $Y=-386400 $D=0
M29 1 IN1 VDD ptft L=1e-05 W=0.0004 $X=10000 $Y=0 $D=0
M30 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=50000 $Y=-386400 $D=0
M31 VDD IN1 1 ptft L=1e-05 W=0.0004 $X=50000 $Y=0 $D=0
M32 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=90000 $Y=-386400 $D=0
M33 1 IN1 VDD ptft L=1e-05 W=0.0004 $X=90000 $Y=0 $D=0
M34 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=130000 $Y=-386400 $D=0
M35 VDD IN1 1 ptft L=1e-05 W=0.0004 $X=130000 $Y=0 $D=0
M36 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=170000 $Y=-386400 $D=0
M37 1 IN1 VDD ptft L=1e-05 W=0.0004 $X=170000 $Y=0 $D=0
M38 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=210000 $Y=-386400 $D=0
M39 VDD IN1 1 ptft L=1e-05 W=0.0004 $X=210000 $Y=0 $D=0
M40 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=250000 $Y=-386400 $D=0
M41 1 IN2 VDD ptft L=1e-05 W=0.0004 $X=250000 $Y=0 $D=0
M42 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=290000 $Y=-386400 $D=0
M43 VDD IN2 1 ptft L=1e-05 W=0.0004 $X=290000 $Y=0 $D=0
M44 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=330000 $Y=-386400 $D=0
M45 1 IN2 VDD ptft L=1e-05 W=0.0004 $X=330000 $Y=0 $D=0
M46 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=370000 $Y=-386400 $D=0
M47 VDD IN2 1 ptft L=1e-05 W=0.0004 $X=370000 $Y=0 $D=0
M48 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=410000 $Y=-386400 $D=0
M49 1 IN2 VDD ptft L=1e-05 W=0.0004 $X=410000 $Y=0 $D=0
M50 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=450000 $Y=-386400 $D=0
M51 VDD IN2 1 ptft L=1e-05 W=0.0004 $X=450000 $Y=0 $D=0
M52 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=490000 $Y=-386400 $D=0
M53 1 IN2 VDD ptft L=1e-05 W=0.0004 $X=490000 $Y=0 $D=0
M54 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=530000 $Y=-386400 $D=0
M55 VDD IN2 1 ptft L=1e-05 W=0.0004 $X=530000 $Y=0 $D=0
M56 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=570000 $Y=-386400 $D=0
M57 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=570000 $Y=0 $D=0
M58 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=610000 $Y=-386400 $D=0
M59 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=610000 $Y=0 $D=0
M60 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=650000 $Y=-386400 $D=0
M61 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=650000 $Y=0 $D=0
M62 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=690000 $Y=-386400 $D=0
M63 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=690000 $Y=0 $D=0
M64 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=730000 $Y=-386400 $D=0
M65 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=730000 $Y=0 $D=0
M66 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=770000 $Y=-386400 $D=0
M67 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=770000 $Y=0 $D=0
M68 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=810000 $Y=-386400 $D=0
M69 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=810000 $Y=0 $D=0
M70 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=850000 $Y=-386400 $D=0
M71 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=850000 $Y=0 $D=0
M72 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=890000 $Y=-386400 $D=0
M73 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=890000 $Y=0 $D=0
M74 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=930000 $Y=-386400 $D=0
M75 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=930000 $Y=0 $D=0
M76 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=970000 $Y=-386400 $D=0
M77 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=970000 $Y=0 $D=0
M78 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1010000 $Y=-386400 $D=0
M79 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=1010000 $Y=0 $D=0
M80 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1050000 $Y=-386400 $D=0
M81 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=1050000 $Y=0 $D=0
M82 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1090000 $Y=-386400 $D=0
M83 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=1090000 $Y=0 $D=0
M84 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1130000 $Y=-386400 $D=0
M85 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=1130000 $Y=0 $D=0
M86 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1170000 $Y=-386400 $D=0
M87 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=1170000 $Y=0 $D=0
.ENDS
***************************************
