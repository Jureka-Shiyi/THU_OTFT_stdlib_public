* File: NAND2D1.cdl
* Created: Sat Aug 17 14:14:15 2024
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "/data/zhengyj/OTFT_stdlib/subckts/NAND2D1.cdl.pex"
.subckt NAND2D1  IN1 IN2 VSS VDD OUT
* 
* OUT	OUT
* VDD	VDD
* VSS	VSS
* IN2	IN2
* IN1	IN1
XMI5 net7 N_IN2_MI5_g N_VSS_MI5_s ntft L=4e-06 W=4e-05
XMI4 N_OUT_MI4_d N_IN1_MI4_g net7 ntft L=4e-06 W=4e-05
XMI2 N_OUT_MI2_d N_IN1_MI2_g N_VDD_MI2_s ptft L=4e-06 W=1e-05
XMI3 N_OUT_MI3_d N_IN2_MI3_g N_VDD_MI3_s ptft L=4e-06 W=1e-05
c_87 net7 0 0.319791f
*
.include "/data/zhengyj/OTFT_stdlib/subckts/NAND2D1.cdl.NAND2D1.pxi"
*
.ends
*
*
