* File: NAND2D4.cdl
* Created: Sat Aug 17 14:17:48 2024
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "/data/zhengyj/OTFT_stdlib/subckts/NAND2D4.cdl.pex"
.subckt NAND2D4  IN1 IN2 VDD OUT VSS
* 
* VSS	VSS
* OUT	OUT
* VDD	VDD
* IN2	IN2
* IN1	IN1
XMI4 N_OUT_MI4_d N_IN1_MI4_g N_net7_MI4_s ntft L=4e-06 W=8e-05
XMI4@2 N_OUT_MI4_d N_IN1_MI4@2_g N_net7_MI4@2_s ntft L=4e-06 W=8e-05
XMI5 N_net7_MI5_d N_IN2_MI5_g N_VSS_MI5_s ntft L=4e-06 W=8e-05
XMI5@2 N_net7_MI5_d N_IN2_MI5@2_g N_VSS_MI5@2_s ntft L=4e-06 W=8e-05
XMI2 N_OUT_MI2_d N_IN1_MI2_g N_VDD_MI2_s ptft L=4e-06 W=4e-05
XMI3 N_OUT_MI3_d N_IN2_MI3_g N_VDD_MI3_s ptft L=4e-06 W=4e-05
*
.include "/data/zhengyj/OTFT_stdlib/subckts/NAND2D4.cdl.NAND2D4.pxi"
*
.ends
*
*
