* SPICE NETLIST
***************************************

.SUBCKT NAND2D4 VSS OUT VDD IN1 IN2
** N=6 EP=5 IP=0 FDC=44
M0 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=-230000 $Y=0 $D=0
M1 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=-190000 $Y=0 $D=0
M2 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=-150000 $Y=0 $D=0
M3 1 VSS VSS ptft L=1e-05 W=0.0001 $X=-144600 $Y=-257600 $D=0
M4 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=-110000 $Y=0 $D=0
M5 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=-104600 $Y=-257600 $D=0
M6 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=-70000 $Y=0 $D=0
M7 1 VSS VSS ptft L=1e-05 W=0.0001 $X=-64600 $Y=-257600 $D=0
M8 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=-30000 $Y=0 $D=0
M9 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=-24600 $Y=-257600 $D=0
M10 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=10000 $Y=0 $D=0
M11 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=50000 $Y=0 $D=0
M12 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=90000 $Y=-386400 $D=0
M13 1 IN1 VDD ptft L=1e-05 W=0.0004 $X=90000 $Y=0 $D=0
M14 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=130000 $Y=-386400 $D=0
M15 VDD IN1 1 ptft L=1e-05 W=0.0004 $X=130000 $Y=0 $D=0
M16 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=170000 $Y=-386400 $D=0
M17 1 IN1 VDD ptft L=1e-05 W=0.0004 $X=170000 $Y=0 $D=0
M18 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=210000 $Y=-386400 $D=0
M19 VDD IN1 1 ptft L=1e-05 W=0.0004 $X=210000 $Y=0 $D=0
M20 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=250000 $Y=-386400 $D=0
M21 1 IN2 VDD ptft L=1e-05 W=0.0004 $X=250000 $Y=0 $D=0
M22 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=290000 $Y=-386400 $D=0
M23 VDD IN2 1 ptft L=1e-05 W=0.0004 $X=290000 $Y=0 $D=0
M24 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=330000 $Y=-386400 $D=0
M25 1 IN2 VDD ptft L=1e-05 W=0.0004 $X=330000 $Y=0 $D=0
M26 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=370000 $Y=-386400 $D=0
M27 VDD IN2 1 ptft L=1e-05 W=0.0004 $X=370000 $Y=0 $D=0
M28 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=410000 $Y=-386400 $D=0
M29 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=410000 $Y=0 $D=0
M30 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=450000 $Y=-386400 $D=0
M31 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=450000 $Y=0 $D=0
M32 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=490000 $Y=-386400 $D=0
M33 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=490000 $Y=0 $D=0
M34 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=530000 $Y=-386400 $D=0
M35 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=530000 $Y=0 $D=0
M36 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=570000 $Y=-386400 $D=0
M37 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=570000 $Y=0 $D=0
M38 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=610000 $Y=-386400 $D=0
M39 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=610000 $Y=0 $D=0
M40 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=650000 $Y=-386400 $D=0
M41 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=650000 $Y=0 $D=0
M42 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=690000 $Y=-386400 $D=0
M43 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=690000 $Y=0 $D=0
.ENDS
***************************************
