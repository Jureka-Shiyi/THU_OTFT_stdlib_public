* SPICE NETLIST
***************************************

.SUBCKT NOR2D2 VSS OUT VDD IN2 IN1
** N=8 EP=5 IP=0 FDC=34
M0 2 VSS VSS ptft L=1e-05 W=0.0002 $X=60000 $Y=160000 $D=0
M1 2 IN2 3 ptft L=1e-05 W=0.0002 $X=70000 $Y=310000 $D=0
M2 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=70000 $Y=630000 $D=0
M3 3 IN2 2 ptft L=1e-05 W=0.0002 $X=110000 $Y=310000 $D=0
M4 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=110000 $Y=630000 $D=0
M5 2 IN2 3 ptft L=1e-05 W=0.0002 $X=150000 $Y=310000 $D=0
M6 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=150000 $Y=630000 $D=0
M7 3 IN2 2 ptft L=1e-05 W=0.0002 $X=190000 $Y=310000 $D=0
M8 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=190000 $Y=630000 $D=0
M9 2 IN2 3 ptft L=1e-05 W=0.0002 $X=230000 $Y=310000 $D=0
M10 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=230000 $Y=630000 $D=0
M11 3 IN2 2 ptft L=1e-05 W=0.0002 $X=270000 $Y=310000 $D=0
M12 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=270000 $Y=630000 $D=0
M13 2 IN2 3 ptft L=1e-05 W=0.0002 $X=310000 $Y=310000 $D=0
M14 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=310000 $Y=630000 $D=0
M15 3 IN2 2 ptft L=1e-05 W=0.0002 $X=350000 $Y=310000 $D=0
M16 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=350000 $Y=630000 $D=0
M17 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=460000 $Y=310000 $D=0
M18 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=460000 $Y=630000 $D=0
M19 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=500000 $Y=310000 $D=0
M20 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=500000 $Y=630000 $D=0
M21 OUT 2 VSS ptft L=1e-05 W=0.0002 $X=525000 $Y=120000 $D=0
M22 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=540000 $Y=310000 $D=0
M23 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=540000 $Y=630000 $D=0
M24 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=580000 $Y=310000 $D=0
M25 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=580000 $Y=630000 $D=0
M26 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=620000 $Y=310000 $D=0
M27 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=620000 $Y=630000 $D=0
M28 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=660000 $Y=310000 $D=0
M29 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=660000 $Y=630000 $D=0
M30 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=700000 $Y=310000 $D=0
M31 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=700000 $Y=630000 $D=0
M32 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=740000 $Y=310000 $D=0
M33 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=740000 $Y=630000 $D=0
.ENDS
***************************************
