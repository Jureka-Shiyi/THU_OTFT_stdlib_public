* File: NAND2D8.cdl
* Created: Mon Dec 22 21:03:44 2025
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "/data/zhengyj/OTFT_stdlib/subckts_cdl/NAND2D8.cdl.pex"
.subckt NAND2D8  VSS OUT VDD IN1 IN2
* 
* IN2	IN2
* IN1	IN1
* VDD	VDD
* OUT	OUT
* VSS	VSS
XMI4 N_OUT_MI4_d N_IN1_MI4_g N_VDD_MI4_s ptft L=1e-05 W=0.0004
XMI4@16 N_OUT_MI4_d N_IN1_MI4@16_g N_VDD_MI4@16_s ptft L=1e-05 W=0.0004
XMI4@15 N_OUT_MI4@15_d N_IN1_MI4@15_g N_VDD_MI4@16_s ptft L=1e-05 W=0.0004
XMI4@14 N_OUT_MI4@15_d N_IN1_MI4@14_g N_VDD_MI4@14_s ptft L=1e-05 W=0.0004
XMI4@13 N_OUT_MI4@13_d N_IN1_MI4@13_g N_VDD_MI4@14_s ptft L=1e-05 W=0.0004
XMI4@12 N_OUT_MI4@13_d N_IN1_MI4@12_g N_VDD_MI4@12_s ptft L=1e-05 W=0.0004
XMI4@11 N_OUT_MI4@11_d N_IN1_MI4@11_g N_VDD_MI4@12_s ptft L=1e-05 W=0.0004
XMI2 N_VSS_MI2_d N_VSS_MI2_g N_net14_MI2_s ptft L=1e-05 W=0.0001
XMI4@10 N_OUT_MI4@11_d N_IN1_MI4@10_g N_VDD_MI4@10_s ptft L=1e-05 W=0.0004
XMI2@8 N_VSS_MI2@8_d N_VSS_MI2@8_g N_net14_MI2_s ptft L=1e-05 W=0.0001
XMI4@9 N_OUT_MI4@9_d N_IN1_MI4@9_g N_VDD_MI4@10_s ptft L=1e-05 W=0.0004
XMI2@7 N_VSS_MI2@8_d N_VSS_MI2@7_g N_net14_MI2@7_s ptft L=1e-05 W=0.0001
XMI4@8 N_OUT_MI4@9_d N_IN1_MI4@8_g N_VDD_MI4@8_s ptft L=1e-05 W=0.0004
XMI2@6 N_VSS_MI2@6_d N_VSS_MI2@6_g N_net14_MI2@7_s ptft L=1e-05 W=0.0001
XMI4@7 N_OUT_MI4@7_d N_IN1_MI4@7_g N_VDD_MI4@8_s ptft L=1e-05 W=0.0004
XMI2@5 N_VSS_MI2@6_d N_VSS_MI2@5_g N_net14_MI2@5_s ptft L=1e-05 W=0.0001
XMI4@6 N_OUT_MI4@7_d N_IN1_MI4@6_g N_VDD_MI4@6_s ptft L=1e-05 W=0.0004
XMI2@4 N_VSS_MI2@4_d N_VSS_MI2@4_g N_net14_MI2@5_s ptft L=1e-05 W=0.0001
XMI4@5 N_OUT_MI4@5_d N_IN1_MI4@5_g N_VDD_MI4@6_s ptft L=1e-05 W=0.0004
XMI2@3 N_VSS_MI2@4_d N_VSS_MI2@3_g N_net14_MI2@3_s ptft L=1e-05 W=0.0001
XMI4@4 N_OUT_MI4@5_d N_IN1_MI4@4_g N_VDD_MI4@4_s ptft L=1e-05 W=0.0004
XMI2@2 N_VSS_MI2@2_d N_VSS_MI2@2_g N_net14_MI2@3_s ptft L=1e-05 W=0.0001
XMI4@3 N_OUT_MI4@3_d N_IN1_MI4@3_g N_VDD_MI4@4_s ptft L=1e-05 W=0.0004
XMI4@2 N_OUT_MI4@3_d N_IN1_MI4@2_g N_VDD_MI4@2_s ptft L=1e-05 W=0.0004
XMI5 N_VSS_MI5_d N_net14_MI5_g N_OUT_MI5_s ptft L=1e-05 W=0.0002
XMI0 N_net14_MI0_d N_IN1_MI0_g N_VDD_MI4@2_s ptft L=1e-05 W=0.0004
XMI5@32 N_VSS_MI5@32_d N_net14_MI5@32_g N_OUT_MI5_s ptft L=1e-05 W=0.0002
XMI0@8 N_net14_MI0_d N_IN1_MI0@8_g N_VDD_MI0@8_s ptft L=1e-05 W=0.0004
XMI5@31 N_VSS_MI5@32_d N_net14_MI5@31_g N_OUT_MI5@31_s ptft L=1e-05 W=0.0002
XMI0@7 N_net14_MI0@7_d N_IN1_MI0@7_g N_VDD_MI0@8_s ptft L=1e-05 W=0.0004
XMI5@30 N_VSS_MI5@30_d N_net14_MI5@30_g N_OUT_MI5@31_s ptft L=1e-05 W=0.0002
XMI0@6 N_net14_MI0@7_d N_IN1_MI0@6_g N_VDD_MI0@6_s ptft L=1e-05 W=0.0004
XMI5@29 N_VSS_MI5@30_d N_net14_MI5@29_g N_OUT_MI5@29_s ptft L=1e-05 W=0.0002
XMI0@5 N_net14_MI0@5_d N_IN1_MI0@5_g N_VDD_MI0@6_s ptft L=1e-05 W=0.0004
XMI5@28 N_VSS_MI5@28_d N_net14_MI5@28_g N_OUT_MI5@29_s ptft L=1e-05 W=0.0002
XMI0@4 N_net14_MI0@5_d N_IN1_MI0@4_g N_VDD_MI0@4_s ptft L=1e-05 W=0.0004
XMI5@27 N_VSS_MI5@28_d N_net14_MI5@27_g N_OUT_MI5@27_s ptft L=1e-05 W=0.0002
XMI0@3 N_net14_MI0@3_d N_IN1_MI0@3_g N_VDD_MI0@4_s ptft L=1e-05 W=0.0004
XMI5@26 N_VSS_MI5@26_d N_net14_MI5@26_g N_OUT_MI5@27_s ptft L=1e-05 W=0.0002
XMI0@2 N_net14_MI0@3_d N_IN1_MI0@2_g N_VDD_MI0@2_s ptft L=1e-05 W=0.0004
XMI5@25 N_VSS_MI5@26_d N_net14_MI5@25_g N_OUT_MI5@25_s ptft L=1e-05 W=0.0002
XMI1 N_net14_MI1_d N_IN2_MI1_g N_VDD_MI0@2_s ptft L=1e-05 W=0.0004
XMI5@24 N_VSS_MI5@24_d N_net14_MI5@24_g N_OUT_MI5@25_s ptft L=1e-05 W=0.0002
XMI1@8 N_net14_MI1_d N_IN2_MI1@8_g N_VDD_MI1@8_s ptft L=1e-05 W=0.0004
XMI5@23 N_VSS_MI5@24_d N_net14_MI5@23_g N_OUT_MI5@23_s ptft L=1e-05 W=0.0002
XMI1@7 N_net14_MI1@7_d N_IN2_MI1@7_g N_VDD_MI1@8_s ptft L=1e-05 W=0.0004
XMI5@22 N_VSS_MI5@22_d N_net14_MI5@22_g N_OUT_MI5@23_s ptft L=1e-05 W=0.0002
XMI1@6 N_net14_MI1@7_d N_IN2_MI1@6_g N_VDD_MI1@6_s ptft L=1e-05 W=0.0004
XMI5@21 N_VSS_MI5@22_d N_net14_MI5@21_g N_OUT_MI5@21_s ptft L=1e-05 W=0.0002
XMI1@5 N_net14_MI1@5_d N_IN2_MI1@5_g N_VDD_MI1@6_s ptft L=1e-05 W=0.0004
XMI5@20 N_VSS_MI5@20_d N_net14_MI5@20_g N_OUT_MI5@21_s ptft L=1e-05 W=0.0002
XMI1@4 N_net14_MI1@5_d N_IN2_MI1@4_g N_VDD_MI1@4_s ptft L=1e-05 W=0.0004
XMI5@19 N_VSS_MI5@20_d N_net14_MI5@19_g N_OUT_MI5@19_s ptft L=1e-05 W=0.0002
XMI1@3 N_net14_MI1@3_d N_IN2_MI1@3_g N_VDD_MI1@4_s ptft L=1e-05 W=0.0004
XMI5@18 N_VSS_MI5@18_d N_net14_MI5@18_g N_OUT_MI5@19_s ptft L=1e-05 W=0.0002
XMI1@2 N_net14_MI1@3_d N_IN2_MI1@2_g N_VDD_MI1@2_s ptft L=1e-05 W=0.0004
XMI5@17 N_VSS_MI5@18_d N_net14_MI5@17_g N_OUT_MI5@17_s ptft L=1e-05 W=0.0002
XMI3 N_OUT_MI3_d N_IN2_MI3_g N_VDD_MI1@2_s ptft L=1e-05 W=0.0004
XMI5@16 N_VSS_MI5@16_d N_net14_MI5@16_g N_OUT_MI5@17_s ptft L=1e-05 W=0.0002
XMI3@16 N_OUT_MI3_d N_IN2_MI3@16_g N_VDD_MI3@16_s ptft L=1e-05 W=0.0004
XMI5@15 N_VSS_MI5@16_d N_net14_MI5@15_g N_OUT_MI5@15_s ptft L=1e-05 W=0.0002
XMI3@15 N_OUT_MI3@15_d N_IN2_MI3@15_g N_VDD_MI3@16_s ptft L=1e-05 W=0.0004
XMI5@14 N_VSS_MI5@14_d N_net14_MI5@14_g N_OUT_MI5@15_s ptft L=1e-05 W=0.0002
XMI3@14 N_OUT_MI3@15_d N_IN2_MI3@14_g N_VDD_MI3@14_s ptft L=1e-05 W=0.0004
XMI5@13 N_VSS_MI5@14_d N_net14_MI5@13_g N_OUT_MI5@13_s ptft L=1e-05 W=0.0002
XMI3@13 N_OUT_MI3@13_d N_IN2_MI3@13_g N_VDD_MI3@14_s ptft L=1e-05 W=0.0004
XMI5@12 N_VSS_MI5@12_d N_net14_MI5@12_g N_OUT_MI5@13_s ptft L=1e-05 W=0.0002
XMI3@12 N_OUT_MI3@13_d N_IN2_MI3@12_g N_VDD_MI3@12_s ptft L=1e-05 W=0.0004
XMI5@11 N_VSS_MI5@12_d N_net14_MI5@11_g N_OUT_MI5@11_s ptft L=1e-05 W=0.0002
XMI3@11 N_OUT_MI3@11_d N_IN2_MI3@11_g N_VDD_MI3@12_s ptft L=1e-05 W=0.0004
XMI5@10 N_VSS_MI5@10_d N_net14_MI5@10_g N_OUT_MI5@11_s ptft L=1e-05 W=0.0002
XMI3@10 N_OUT_MI3@11_d N_IN2_MI3@10_g N_VDD_MI3@10_s ptft L=1e-05 W=0.0004
XMI5@9 N_VSS_MI5@10_d N_net14_MI5@9_g N_OUT_MI5@9_s ptft L=1e-05 W=0.0002
XMI3@9 N_OUT_MI3@9_d N_IN2_MI3@9_g N_VDD_MI3@10_s ptft L=1e-05 W=0.0004
XMI5@8 N_VSS_MI5@8_d N_net14_MI5@8_g N_OUT_MI5@9_s ptft L=1e-05 W=0.0002
XMI3@8 N_OUT_MI3@9_d N_IN2_MI3@8_g N_VDD_MI3@8_s ptft L=1e-05 W=0.0004
XMI5@7 N_VSS_MI5@8_d N_net14_MI5@7_g N_OUT_MI5@7_s ptft L=1e-05 W=0.0002
XMI3@7 N_OUT_MI3@7_d N_IN2_MI3@7_g N_VDD_MI3@8_s ptft L=1e-05 W=0.0004
XMI5@6 N_VSS_MI5@6_d N_net14_MI5@6_g N_OUT_MI5@7_s ptft L=1e-05 W=0.0002
XMI3@6 N_OUT_MI3@7_d N_IN2_MI3@6_g N_VDD_MI3@6_s ptft L=1e-05 W=0.0004
XMI5@5 N_VSS_MI5@6_d N_net14_MI5@5_g N_OUT_MI5@5_s ptft L=1e-05 W=0.0002
XMI3@5 N_OUT_MI3@5_d N_IN2_MI3@5_g N_VDD_MI3@6_s ptft L=1e-05 W=0.0004
XMI5@4 N_VSS_MI5@4_d N_net14_MI5@4_g N_OUT_MI5@5_s ptft L=1e-05 W=0.0002
XMI3@4 N_OUT_MI3@5_d N_IN2_MI3@4_g N_VDD_MI3@4_s ptft L=1e-05 W=0.0004
XMI5@3 N_VSS_MI5@4_d N_net14_MI5@3_g N_OUT_MI5@3_s ptft L=1e-05 W=0.0002
XMI3@3 N_OUT_MI3@3_d N_IN2_MI3@3_g N_VDD_MI3@4_s ptft L=1e-05 W=0.0004
XMI5@2 N_VSS_MI5@2_d N_net14_MI5@2_g N_OUT_MI5@3_s ptft L=1e-05 W=0.0002
XMI3@2 N_OUT_MI3@3_d N_IN2_MI3@2_g N_VDD_MI3@2_s ptft L=1e-05 W=0.0004
*
.include "/data/zhengyj/OTFT_stdlib/subckts_cdl/NAND2D8.cdl.NAND2D8.pxi"
*
.ends
*
*
