* File: NOR2D8.cdl
* Created: Mon Dec 22 21:23:22 2025
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "/data/zhengyj/OTFT_stdlib/subckts_cdl/NOR2D8.cdl.pex"
.subckt NOR2D8  VSS OUT VDD IN2 IN1
* 
* IN1	IN1
* IN2	IN2
* VDD	VDD
* OUT	OUT
* VSS	VSS
XMI4 N_VSS_MI4_d N_VSS_MI4_g N_net11_MI4_s ptft L=1e-05 W=0.0008
XMI1 N_net11_MI1_d N_IN2_MI1_g N_net10_MI1_s ptft L=1e-05 W=0.0002
XMI0 N_net10_MI0_d N_IN1_MI0_g N_VDD_MI0_s ptft L=1e-05 W=0.0002
XMI1@32 N_net11_MI1_d N_IN2_MI1@32_g N_net10_MI1@32_s ptft L=1e-05 W=0.0002
XMI0@32 N_net10_MI0@32_d N_IN1_MI0@32_g N_VDD_MI0_s ptft L=1e-05 W=0.0002
XMI1@31 N_net11_MI1@31_d N_IN2_MI1@31_g N_net10_MI1@32_s ptft L=1e-05 W=0.0002
XMI0@31 N_net10_MI0@32_d N_IN1_MI0@31_g N_VDD_MI0@31_s ptft L=1e-05 W=0.0002
XMI1@30 N_net11_MI1@31_d N_IN2_MI1@30_g N_net10_MI1@30_s ptft L=1e-05 W=0.0002
XMI0@30 N_net10_MI0@30_d N_IN1_MI0@30_g N_VDD_MI0@31_s ptft L=1e-05 W=0.0002
XMI1@29 N_net11_MI1@29_d N_IN2_MI1@29_g N_net10_MI1@30_s ptft L=1e-05 W=0.0002
XMI0@29 N_net10_MI0@30_d N_IN1_MI0@29_g N_VDD_MI0@29_s ptft L=1e-05 W=0.0002
XMI1@28 N_net11_MI1@29_d N_IN2_MI1@28_g N_net10_MI1@28_s ptft L=1e-05 W=0.0002
XMI0@28 N_net10_MI0@28_d N_IN1_MI0@28_g N_VDD_MI0@29_s ptft L=1e-05 W=0.0002
XMI1@27 N_net11_MI1@27_d N_IN2_MI1@27_g N_net10_MI1@28_s ptft L=1e-05 W=0.0002
XMI0@27 N_net10_MI0@28_d N_IN1_MI0@27_g N_VDD_MI0@27_s ptft L=1e-05 W=0.0002
XMI1@26 N_net11_MI1@27_d N_IN2_MI1@26_g N_net10_MI1@26_s ptft L=1e-05 W=0.0002
XMI0@26 N_net10_MI0@26_d N_IN1_MI0@26_g N_VDD_MI0@27_s ptft L=1e-05 W=0.0002
XMI1@25 N_net11_MI1@25_d N_IN2_MI1@25_g N_net10_MI1@26_s ptft L=1e-05 W=0.0002
XMI0@25 N_net10_MI0@26_d N_IN1_MI0@25_g N_VDD_MI0@25_s ptft L=1e-05 W=0.0002
XMI1@24 N_net11_MI1@25_d N_IN2_MI1@24_g N_net10_MI1@24_s ptft L=1e-05 W=0.0002
XMI0@24 N_net10_MI0@24_d N_IN1_MI0@24_g N_VDD_MI0@25_s ptft L=1e-05 W=0.0002
XMI1@23 N_net11_MI1@23_d N_IN2_MI1@23_g N_net10_MI1@24_s ptft L=1e-05 W=0.0002
XMI0@23 N_net10_MI0@24_d N_IN1_MI0@23_g N_VDD_MI0@23_s ptft L=1e-05 W=0.0002
XMI1@22 N_net11_MI1@23_d N_IN2_MI1@22_g N_net10_MI1@22_s ptft L=1e-05 W=0.0002
XMI0@22 N_net10_MI0@22_d N_IN1_MI0@22_g N_VDD_MI0@23_s ptft L=1e-05 W=0.0002
XMI1@21 N_net11_MI1@21_d N_IN2_MI1@21_g N_net10_MI1@22_s ptft L=1e-05 W=0.0002
XMI0@21 N_net10_MI0@22_d N_IN1_MI0@21_g N_VDD_MI0@21_s ptft L=1e-05 W=0.0002
XMI1@20 N_net11_MI1@21_d N_IN2_MI1@20_g N_net10_MI1@20_s ptft L=1e-05 W=0.0002
XMI0@20 N_net10_MI0@20_d N_IN1_MI0@20_g N_VDD_MI0@21_s ptft L=1e-05 W=0.0002
XMI1@19 N_net11_MI1@19_d N_IN2_MI1@19_g N_net10_MI1@20_s ptft L=1e-05 W=0.0002
XMI0@19 N_net10_MI0@20_d N_IN1_MI0@19_g N_VDD_MI0@19_s ptft L=1e-05 W=0.0002
XMI1@18 N_net11_MI1@19_d N_IN2_MI1@18_g N_net10_MI1@18_s ptft L=1e-05 W=0.0002
XMI0@18 N_net10_MI0@18_d N_IN1_MI0@18_g N_VDD_MI0@19_s ptft L=1e-05 W=0.0002
XMI1@17 N_net11_MI1@17_d N_IN2_MI1@17_g N_net10_MI1@18_s ptft L=1e-05 W=0.0002
XMI0@17 N_net10_MI0@18_d N_IN1_MI0@17_g N_VDD_MI0@17_s ptft L=1e-05 W=0.0002
XMI1@16 N_net11_MI1@17_d N_IN2_MI1@16_g N_net10_MI1@16_s ptft L=1e-05 W=0.0002
XMI0@16 N_net10_MI0@16_d N_IN1_MI0@16_g N_VDD_MI0@17_s ptft L=1e-05 W=0.0002
XMI1@15 N_net11_MI1@15_d N_IN2_MI1@15_g N_net10_MI1@16_s ptft L=1e-05 W=0.0002
XMI0@15 N_net10_MI0@16_d N_IN1_MI0@15_g N_VDD_MI0@15_s ptft L=1e-05 W=0.0002
XMI1@14 N_net11_MI1@15_d N_IN2_MI1@14_g N_net10_MI1@14_s ptft L=1e-05 W=0.0002
XMI0@14 N_net10_MI0@14_d N_IN1_MI0@14_g N_VDD_MI0@15_s ptft L=1e-05 W=0.0002
XMI1@13 N_net11_MI1@13_d N_IN2_MI1@13_g N_net10_MI1@14_s ptft L=1e-05 W=0.0002
XMI0@13 N_net10_MI0@14_d N_IN1_MI0@13_g N_VDD_MI0@13_s ptft L=1e-05 W=0.0002
XMI1@12 N_net11_MI1@13_d N_IN2_MI1@12_g N_net10_MI1@12_s ptft L=1e-05 W=0.0002
XMI0@12 N_net10_MI0@12_d N_IN1_MI0@12_g N_VDD_MI0@13_s ptft L=1e-05 W=0.0002
XMI1@11 N_net11_MI1@11_d N_IN2_MI1@11_g N_net10_MI1@12_s ptft L=1e-05 W=0.0002
XMI0@11 N_net10_MI0@12_d N_IN1_MI0@11_g N_VDD_MI0@11_s ptft L=1e-05 W=0.0002
XMI1@10 N_net11_MI1@11_d N_IN2_MI1@10_g N_net10_MI1@10_s ptft L=1e-05 W=0.0002
XMI0@10 N_net10_MI0@10_d N_IN1_MI0@10_g N_VDD_MI0@11_s ptft L=1e-05 W=0.0002
XMI1@9 N_net11_MI1@9_d N_IN2_MI1@9_g N_net10_MI1@10_s ptft L=1e-05 W=0.0002
XMI0@9 N_net10_MI0@10_d N_IN1_MI0@9_g N_VDD_MI0@9_s ptft L=1e-05 W=0.0002
XMI1@8 N_net11_MI1@9_d N_IN2_MI1@8_g N_net10_MI1@8_s ptft L=1e-05 W=0.0002
XMI0@8 N_net10_MI0@8_d N_IN1_MI0@8_g N_VDD_MI0@9_s ptft L=1e-05 W=0.0002
XMI1@7 N_net11_MI1@7_d N_IN2_MI1@7_g N_net10_MI1@8_s ptft L=1e-05 W=0.0002
XMI0@7 N_net10_MI0@8_d N_IN1_MI0@7_g N_VDD_MI0@7_s ptft L=1e-05 W=0.0002
XMI1@6 N_net11_MI1@7_d N_IN2_MI1@6_g N_net10_MI1@6_s ptft L=1e-05 W=0.0002
XMI0@6 N_net10_MI0@6_d N_IN1_MI0@6_g N_VDD_MI0@7_s ptft L=1e-05 W=0.0002
XMI1@5 N_net11_MI1@5_d N_IN2_MI1@5_g N_net10_MI1@6_s ptft L=1e-05 W=0.0002
XMI0@5 N_net10_MI0@6_d N_IN1_MI0@5_g N_VDD_MI0@5_s ptft L=1e-05 W=0.0002
XMI1@4 N_net11_MI1@5_d N_IN2_MI1@4_g N_net10_MI1@4_s ptft L=1e-05 W=0.0002
XMI0@4 N_net10_MI0@4_d N_IN1_MI0@4_g N_VDD_MI0@5_s ptft L=1e-05 W=0.0002
XMI1@3 N_net11_MI1@3_d N_IN2_MI1@3_g N_net10_MI1@4_s ptft L=1e-05 W=0.0002
XMI0@3 N_net10_MI0@4_d N_IN1_MI0@3_g N_VDD_MI0@3_s ptft L=1e-05 W=0.0002
XMI1@2 N_net11_MI1@3_d N_IN2_MI1@2_g N_net10_MI1@2_s ptft L=1e-05 W=0.0002
XMI0@2 N_net10_MI0@2_d N_IN1_MI0@2_g N_VDD_MI0@3_s ptft L=1e-05 W=0.0002
XMI3 N_OUT_MI3_d N_IN2_MI3_g N_net12_MI3_s ptft L=1e-05 W=0.0002
XMI2 N_net12_MI2_d N_IN1_MI2_g N_VDD_MI2_s ptft L=1e-05 W=0.0002
XMI3@32 N_OUT_MI3_d N_IN2_MI3@32_g N_net12_MI3@32_s ptft L=1e-05 W=0.0002
XMI2@32 N_net12_MI2@32_d N_IN1_MI2@32_g N_VDD_MI2_s ptft L=1e-05 W=0.0002
XMI3@31 N_OUT_MI3@31_d N_IN2_MI3@31_g N_net12_MI3@32_s ptft L=1e-05 W=0.0002
XMI2@31 N_net12_MI2@32_d N_IN1_MI2@31_g N_VDD_MI2@31_s ptft L=1e-05 W=0.0002
XMI3@30 N_OUT_MI3@31_d N_IN2_MI3@30_g N_net12_MI3@30_s ptft L=1e-05 W=0.0002
XMI2@30 N_net12_MI2@30_d N_IN1_MI2@30_g N_VDD_MI2@31_s ptft L=1e-05 W=0.0002
XMI3@29 N_OUT_MI3@29_d N_IN2_MI3@29_g N_net12_MI3@30_s ptft L=1e-05 W=0.0002
XMI2@29 N_net12_MI2@30_d N_IN1_MI2@29_g N_VDD_MI2@29_s ptft L=1e-05 W=0.0002
XMI3@28 N_OUT_MI3@29_d N_IN2_MI3@28_g N_net12_MI3@28_s ptft L=1e-05 W=0.0002
XMI2@28 N_net12_MI2@28_d N_IN1_MI2@28_g N_VDD_MI2@29_s ptft L=1e-05 W=0.0002
XMI3@27 N_OUT_MI3@27_d N_IN2_MI3@27_g N_net12_MI3@28_s ptft L=1e-05 W=0.0002
XMI2@27 N_net12_MI2@28_d N_IN1_MI2@27_g N_VDD_MI2@27_s ptft L=1e-05 W=0.0002
XMI5 N_VSS_MI5_d N_net11_MI5_g N_OUT_MI5_s ptft L=1e-05 W=0.0008
XMI3@26 N_OUT_MI3@27_d N_IN2_MI3@26_g N_net12_MI3@26_s ptft L=1e-05 W=0.0002
XMI2@26 N_net12_MI2@26_d N_IN1_MI2@26_g N_VDD_MI2@27_s ptft L=1e-05 W=0.0002
XMI3@25 N_OUT_MI3@25_d N_IN2_MI3@25_g N_net12_MI3@26_s ptft L=1e-05 W=0.0002
XMI2@25 N_net12_MI2@26_d N_IN1_MI2@25_g N_VDD_MI2@25_s ptft L=1e-05 W=0.0002
XMI3@24 N_OUT_MI3@25_d N_IN2_MI3@24_g N_net12_MI3@24_s ptft L=1e-05 W=0.0002
XMI2@24 N_net12_MI2@24_d N_IN1_MI2@24_g N_VDD_MI2@25_s ptft L=1e-05 W=0.0002
XMI3@23 N_OUT_MI3@23_d N_IN2_MI3@23_g N_net12_MI3@24_s ptft L=1e-05 W=0.0002
XMI2@23 N_net12_MI2@24_d N_IN1_MI2@23_g N_VDD_MI2@23_s ptft L=1e-05 W=0.0002
XMI3@22 N_OUT_MI3@23_d N_IN2_MI3@22_g N_net12_MI3@22_s ptft L=1e-05 W=0.0002
XMI2@22 N_net12_MI2@22_d N_IN1_MI2@22_g N_VDD_MI2@23_s ptft L=1e-05 W=0.0002
XMI3@21 N_OUT_MI3@21_d N_IN2_MI3@21_g N_net12_MI3@22_s ptft L=1e-05 W=0.0002
XMI2@21 N_net12_MI2@22_d N_IN1_MI2@21_g N_VDD_MI2@21_s ptft L=1e-05 W=0.0002
XMI3@20 N_OUT_MI3@21_d N_IN2_MI3@20_g N_net12_MI3@20_s ptft L=1e-05 W=0.0002
XMI2@20 N_net12_MI2@20_d N_IN1_MI2@20_g N_VDD_MI2@21_s ptft L=1e-05 W=0.0002
XMI3@19 N_OUT_MI3@19_d N_IN2_MI3@19_g N_net12_MI3@20_s ptft L=1e-05 W=0.0002
XMI2@19 N_net12_MI2@20_d N_IN1_MI2@19_g N_VDD_MI2@19_s ptft L=1e-05 W=0.0002
XMI3@18 N_OUT_MI3@19_d N_IN2_MI3@18_g N_net12_MI3@18_s ptft L=1e-05 W=0.0002
XMI2@18 N_net12_MI2@18_d N_IN1_MI2@18_g N_VDD_MI2@19_s ptft L=1e-05 W=0.0002
XMI3@17 N_OUT_MI3@17_d N_IN2_MI3@17_g N_net12_MI3@18_s ptft L=1e-05 W=0.0002
XMI2@17 N_net12_MI2@18_d N_IN1_MI2@17_g N_VDD_MI2@17_s ptft L=1e-05 W=0.0002
XMI3@16 N_OUT_MI3@17_d N_IN2_MI3@16_g N_net12_MI3@16_s ptft L=1e-05 W=0.0002
XMI2@16 N_net12_MI2@16_d N_IN1_MI2@16_g N_VDD_MI2@17_s ptft L=1e-05 W=0.0002
XMI3@15 N_OUT_MI3@15_d N_IN2_MI3@15_g N_net12_MI3@16_s ptft L=1e-05 W=0.0002
XMI2@15 N_net12_MI2@16_d N_IN1_MI2@15_g N_VDD_MI2@15_s ptft L=1e-05 W=0.0002
XMI3@14 N_OUT_MI3@15_d N_IN2_MI3@14_g N_net12_MI3@14_s ptft L=1e-05 W=0.0002
XMI2@14 N_net12_MI2@14_d N_IN1_MI2@14_g N_VDD_MI2@15_s ptft L=1e-05 W=0.0002
XMI3@13 N_OUT_MI3@13_d N_IN2_MI3@13_g N_net12_MI3@14_s ptft L=1e-05 W=0.0002
XMI2@13 N_net12_MI2@14_d N_IN1_MI2@13_g N_VDD_MI2@13_s ptft L=1e-05 W=0.0002
XMI3@12 N_OUT_MI3@13_d N_IN2_MI3@12_g N_net12_MI3@12_s ptft L=1e-05 W=0.0002
XMI2@12 N_net12_MI2@12_d N_IN1_MI2@12_g N_VDD_MI2@13_s ptft L=1e-05 W=0.0002
XMI3@11 N_OUT_MI3@11_d N_IN2_MI3@11_g N_net12_MI3@12_s ptft L=1e-05 W=0.0002
XMI2@11 N_net12_MI2@12_d N_IN1_MI2@11_g N_VDD_MI2@11_s ptft L=1e-05 W=0.0002
XMI3@10 N_OUT_MI3@11_d N_IN2_MI3@10_g N_net12_MI3@10_s ptft L=1e-05 W=0.0002
XMI2@10 N_net12_MI2@10_d N_IN1_MI2@10_g N_VDD_MI2@11_s ptft L=1e-05 W=0.0002
XMI3@9 N_OUT_MI3@9_d N_IN2_MI3@9_g N_net12_MI3@10_s ptft L=1e-05 W=0.0002
XMI2@9 N_net12_MI2@10_d N_IN1_MI2@9_g N_VDD_MI2@9_s ptft L=1e-05 W=0.0002
XMI3@8 N_OUT_MI3@9_d N_IN2_MI3@8_g N_net12_MI3@8_s ptft L=1e-05 W=0.0002
XMI2@8 N_net12_MI2@8_d N_IN1_MI2@8_g N_VDD_MI2@9_s ptft L=1e-05 W=0.0002
XMI3@7 N_OUT_MI3@7_d N_IN2_MI3@7_g N_net12_MI3@8_s ptft L=1e-05 W=0.0002
XMI2@7 N_net12_MI2@8_d N_IN1_MI2@7_g N_VDD_MI2@7_s ptft L=1e-05 W=0.0002
XMI3@6 N_OUT_MI3@7_d N_IN2_MI3@6_g N_net12_MI3@6_s ptft L=1e-05 W=0.0002
XMI2@6 N_net12_MI2@6_d N_IN1_MI2@6_g N_VDD_MI2@7_s ptft L=1e-05 W=0.0002
XMI3@5 N_OUT_MI3@5_d N_IN2_MI3@5_g N_net12_MI3@6_s ptft L=1e-05 W=0.0002
XMI2@5 N_net12_MI2@6_d N_IN1_MI2@5_g N_VDD_MI2@5_s ptft L=1e-05 W=0.0002
XMI3@4 N_OUT_MI3@5_d N_IN2_MI3@4_g N_net12_MI3@4_s ptft L=1e-05 W=0.0002
XMI2@4 N_net12_MI2@4_d N_IN1_MI2@4_g N_VDD_MI2@5_s ptft L=1e-05 W=0.0002
XMI3@3 N_OUT_MI3@3_d N_IN2_MI3@3_g N_net12_MI3@4_s ptft L=1e-05 W=0.0002
XMI2@3 N_net12_MI2@4_d N_IN1_MI2@3_g N_VDD_MI2@3_s ptft L=1e-05 W=0.0002
XMI3@2 N_OUT_MI3@3_d N_IN2_MI3@2_g N_net12_MI3@2_s ptft L=1e-05 W=0.0002
XMI2@2 N_net12_MI2@2_d N_IN1_MI2@2_g N_VDD_MI2@3_s ptft L=1e-05 W=0.0002
*
.include "/data/zhengyj/OTFT_stdlib/subckts_cdl/NOR2D8.cdl.NOR2D8.pxi"
*
.ends
*
*
