* File: XOR2D8.cdl
* Created: Thu Jan 16 00:33:32 2025
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "/data/zhengyj/OTFT_stdlib/subckts/XOR2D8.cdl.pex"
.subckt XOR2D8  IN2 IN1 VSS VDD OUT
* 
* OUT	OUT
* VDD	VDD
* VSS	VSS
* IN1	IN1
* IN2	IN2
XMI5 N_net23_MI5_d N_IN1_MI5_g N_VSS_MI5_s ntft L=4e-06 W=8e-05
XMI1 N_net23_MI1_d N_IN1_MI1_g N_VSS_MI1_s ntft L=4e-06 W=8e-05
XMI16 N_net25_MI16_d N_IN2_MI16_g N_VSS_MI16_s ntft L=4e-06 W=8e-05
XMI15 N_net25_MI15_d N_IN2_MI15_g N_VSS_MI15_s ntft L=4e-06 W=8e-05
XMI23 N_net23_MI23_d N_net25_MI23_g N_net26_MI23_s ntft L=4e-06 W=8e-05
XMI11 N_net23_MI11_d N_net25_MI11_g N_net26_MI11_s ntft L=4e-06 W=8e-05
XMI26 N_OUT_MI26_d N_net26_MI26_g N_VSS_MI26_s ntft L=4e-06 W=8e-05
XMI25 N_OUT_MI25_d N_net26_MI25_g N_VSS_MI25_s ntft L=4e-06 W=8e-05
XMI13 N_OUT_MI13_d N_net26_MI13_g N_VSS_MI13_s ntft L=4e-06 W=8e-05
XMI4 N_OUT_MI4_d N_net26_MI4_g N_VSS_MI4_s ntft L=4e-06 W=8e-05
XMI0 N_net23_MI0_d N_IN1_MI0_g N_VDD_MI0_s ptft L=4e-06 W=8e-05
XMI14 N_net25_MI14_d N_IN2_MI14_g N_VDD_MI14_s ptft L=4e-06 W=8e-05
XMI18 N_net26_MI18_d N_net25_MI18_g N_net24_MI18_s ptft L=4e-06 W=8e-05
XMI17 N_net24_MI18_s N_net23_MI17_g N_VDD_MI17_s ptft L=4e-06 W=8e-05
XMI7 N_net26_MI7_d N_net25_MI7_g N_net24_MI7_s ptft L=4e-06 W=8e-05
XMI6 N_net24_MI7_s N_net23_MI6_g N_VDD_MI6_s ptft L=4e-06 W=8e-05
XMI10 N_net23_MI10_d N_IN2_MI10_g N_net26_MI10_s ptft L=4e-06 W=8e-05
XMI24 N_OUT_MI24_d N_net26_MI24_g N_VDD_MI24_s ptft L=4e-06 W=8e-05
XMI12 N_OUT_MI12_d N_net26_MI12_g N_VDD_MI12_s ptft L=4e-06 W=8e-05
XMI22 N_net27_MI22_d N_net23_MI22_g N_VSS_MI22_s ntft L=4e-06 W=8e-05
XMI20 N_net26_MI20_d N_IN2_MI20_g N_net27_MI22_d ntft L=4e-06 W=8e-05
XMI21 N_net27_MI21_d N_net23_MI21_g N_VSS_MI21_s ntft L=4e-06 W=8e-05
XMI19 N_net26_MI19_d N_IN2_MI19_g N_net27_MI21_d ntft L=4e-06 W=8e-05
XMI9 N_net27_MI9_d N_net23_MI9_g N_VSS_MI9_s ntft L=4e-06 W=8e-05
XMI8 N_net26_MI8_d N_IN2_MI8_g N_net27_MI9_d ntft L=4e-06 W=8e-05
XMI3 N_net27_MI3_d N_net23_MI3_g N_VSS_MI3_s ntft L=4e-06 W=8e-05
XMI2 N_net26_MI2_d N_IN2_MI2_g N_net27_MI3_d ntft L=4e-06 W=8e-05
*
.include "/data/zhengyj/OTFT_stdlib/subckts/XOR2D8.cdl.XOR2D8.pxi"
*
.ends
*
*
