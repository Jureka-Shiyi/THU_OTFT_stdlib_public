* SPICE NETLIST
***************************************

.SUBCKT BUFD4 VSS VDD OUT IN
** N=7 EP=4 IP=0 FDC=48
M0 1 VSS VSS ptft L=4e-05 W=0.0001 $X=68000 $Y=300000 $D=0
M1 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=148000 $Y=300000 $D=0
M2 VDD IN 1 ptft L=1e-05 W=0.0002 $X=158000 $Y=580000 $D=0
M3 1 IN VDD ptft L=1e-05 W=0.0002 $X=208000 $Y=580000 $D=0
M4 1 VSS VSS ptft L=4e-05 W=0.0001 $X=228000 $Y=300000 $D=0
M5 VDD IN 1 ptft L=1e-05 W=0.0002 $X=258000 $Y=580000 $D=0
M6 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=308000 $Y=300000 $D=0
M7 1 IN VDD ptft L=1e-05 W=0.0002 $X=308000 $Y=580000 $D=0
M8 VSS 1 3 ptft L=1e-05 W=0.0002 $X=478000 $Y=180000 $D=0
M9 VDD IN 3 ptft L=1e-05 W=0.0002 $X=478000 $Y=580000 $D=0
M10 3 1 VSS ptft L=1e-05 W=0.0002 $X=528000 $Y=180000 $D=0
M11 3 IN VDD ptft L=1e-05 W=0.0002 $X=528000 $Y=580000 $D=0
M12 VSS 1 3 ptft L=1e-05 W=0.0002 $X=578000 $Y=180000 $D=0
M13 VDD IN 3 ptft L=1e-05 W=0.0002 $X=578000 $Y=580000 $D=0
M14 3 1 VSS ptft L=1e-05 W=0.0002 $X=628000 $Y=180000 $D=0
M15 3 IN VDD ptft L=1e-05 W=0.0002 $X=628000 $Y=580000 $D=0
M16 VSS 1 3 ptft L=1e-05 W=0.0002 $X=678000 $Y=180000 $D=0
M17 VDD IN 3 ptft L=1e-05 W=0.0002 $X=678000 $Y=580000 $D=0
M18 3 1 VSS ptft L=1e-05 W=0.0002 $X=728000 $Y=180000 $D=0
M19 3 IN VDD ptft L=1e-05 W=0.0002 $X=728000 $Y=580000 $D=0
M20 VSS 1 3 ptft L=1e-05 W=0.0002 $X=778000 $Y=180000 $D=0
M21 VDD IN 3 ptft L=1e-05 W=0.0002 $X=778000 $Y=580000 $D=0
M22 3 1 VSS ptft L=1e-05 W=0.0002 $X=828000 $Y=180000 $D=0
M23 3 IN VDD ptft L=1e-05 W=0.0002 $X=828000 $Y=580000 $D=0
M24 4 VSS VSS ptft L=4e-05 W=0.0001 $X=976000 $Y=300000 $D=0
M25 VSS VSS 4 ptft L=4e-05 W=0.0001 $X=1056000 $Y=300000 $D=0
M26 VDD 3 4 ptft L=1e-05 W=0.0002 $X=1066000 $Y=580000 $D=0
M27 4 3 VDD ptft L=1e-05 W=0.0002 $X=1116000 $Y=580000 $D=0
M28 4 VSS VSS ptft L=4e-05 W=0.0001 $X=1136000 $Y=300000 $D=0
M29 VDD 3 4 ptft L=1e-05 W=0.0002 $X=1166000 $Y=580000 $D=0
M30 VSS VSS 4 ptft L=4e-05 W=0.0001 $X=1216000 $Y=300000 $D=0
M31 4 3 VDD ptft L=1e-05 W=0.0002 $X=1216000 $Y=580000 $D=0
M32 VSS 4 OUT ptft L=1e-05 W=0.0002 $X=1386000 $Y=180000 $D=0
M33 VDD 3 OUT ptft L=1e-05 W=0.0002 $X=1386000 $Y=580000 $D=0
M34 OUT 4 VSS ptft L=1e-05 W=0.0002 $X=1436000 $Y=180000 $D=0
M35 OUT 3 VDD ptft L=1e-05 W=0.0002 $X=1436000 $Y=580000 $D=0
M36 VSS 4 OUT ptft L=1e-05 W=0.0002 $X=1486000 $Y=180000 $D=0
M37 VDD 3 OUT ptft L=1e-05 W=0.0002 $X=1486000 $Y=580000 $D=0
M38 OUT 4 VSS ptft L=1e-05 W=0.0002 $X=1536000 $Y=180000 $D=0
M39 OUT 3 VDD ptft L=1e-05 W=0.0002 $X=1536000 $Y=580000 $D=0
M40 VSS 4 OUT ptft L=1e-05 W=0.0002 $X=1586000 $Y=180000 $D=0
M41 VDD 3 OUT ptft L=1e-05 W=0.0002 $X=1586000 $Y=580000 $D=0
M42 OUT 4 VSS ptft L=1e-05 W=0.0002 $X=1636000 $Y=180000 $D=0
M43 OUT 3 VDD ptft L=1e-05 W=0.0002 $X=1636000 $Y=580000 $D=0
M44 VSS 4 OUT ptft L=1e-05 W=0.0002 $X=1686000 $Y=180000 $D=0
M45 VDD 3 OUT ptft L=1e-05 W=0.0002 $X=1686000 $Y=580000 $D=0
M46 OUT 4 VSS ptft L=1e-05 W=0.0002 $X=1736000 $Y=180000 $D=0
M47 OUT 3 VDD ptft L=1e-05 W=0.0002 $X=1736000 $Y=580000 $D=0
.ENDS
***************************************
