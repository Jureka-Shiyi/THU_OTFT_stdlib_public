* File: DFFD1.cdl
* Created: Sat Dec 27 12:52:46 2025
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "DFFD1.cdl.pex"
.subckt DFFD1  CK D VSS VDD QN Q
* 
* Q	Q
* QN	QN
* VDD	VDD
* VSS	VSS
* D	D
* CK	CK
XMI44 N_net156_MI44_d N_:CK_MI44_g N_VDD_MI44_s ptft L=1.8e-05 W=0.00016
XMI22 N_net167_MI22_d N_CK_MI22_g N_VDD_MI22_s ptft L=1.8e-05 W=0.00016
XMI4 N_net169_MI4_d N_D_MI4_g N_VDD_MI4_s ptft L=1.8e-05 W=0.00016
XMI42 N_VSS_MI42_d N_VSS_MI42_g N_net156_MI42_s ptft L=1.8e-05 W=4e-05
XMI20 N_VSS_MI20_d N_VSS_MI20_g N_net167_MI20_s ptft L=1.8e-05 W=4e-05
XMI5 N_VSS_MI5_d N_VSS_MI5_g N_net169_MI5_s ptft L=1.8e-05 W=4e-05
XMI43 N_VSS_MI43_d N_net156_MI43_g N_::CK_MI43_s ptft L=1.8e-05 W=0.00032
XMI45 N_::CK_MI43_s N_:CK_MI45_g N_VDD_MI45_s ptft L=1.8e-05 W=0.00032
XMI21 N_VSS_MI21_d N_net167_MI21_g N_:CK_MI21_s ptft L=1.8e-05 W=0.00032
XMI23 N_:CK_MI21_s N_CK_MI23_g N_VDD_MI23_s ptft L=1.8e-05 W=0.00032
XMI7 N_VSS_MI7_d N_net169_MI7_g N_:D_MI7_s ptft L=1.8e-05 W=0.00032
XMI6 N_:D_MI7_s N_D_MI6_g N_VDD_MI6_s ptft L=1.8e-05 W=0.00032
XMI27 N_net168_MI27_d N_:CK_MI27_g N_VDD_MI27_s ptft L=1.8e-05 W=0.00012
XMI3 N_net170_MI3_d N_:CK_MI3_g N_VDD_MI3_s ptft L=1.8e-05 W=0.00012
XMI24 N_VSS_MI24_d N_VSS_MI24_g N_net168_MI24_s ptft L=1.8e-05 W=4e-05
XMI2 N_VSS_MI24_d N_VSS_MI2_g N_net170_MI2_s ptft L=1.8e-05 W=4e-05
XMI26 N_net168_MI26_d N_:D_MI26_g N_VDD_MI26_s ptft L=1.8e-05 W=0.00012
XMI1 N_net170_MI1_d N_D_MI1_g N_VDD_MI1_s ptft L=1.8e-05 W=0.00012
XMI29 N_F1N_MI29_d N_:D_MI29_g N_VDD_MI29_s ptft L=1.8e-05 W=0.00024
XMI9 N_F1_MI9_d N_D_MI9_g N_VDD_MI9_s ptft L=1.8e-05 W=0.00024
XMI25 N_VSS_MI25_d N_net168_MI25_g N_F1N_MI25_s ptft L=1.8e-05 W=0.00048
XMI0 N_VSS_MI25_d N_net170_MI0_g N_F1_MI0_s ptft L=1.8e-05 W=0.00048
XMI28 N_F1N_MI28_d N_:CK_MI28_g N_VDD_MI28_s ptft L=1.8e-05 W=0.00024
XMI8 N_F1_MI8_d N_:CK_MI8_g N_VDD_MI8_s ptft L=1.8e-05 W=0.00024
XMI38 N_net160_MI38_d N_F1O_MI38_g N_VDD_MI38_s ptft L=1.8e-05 W=0.00012
XMI33 N_net159_MI33_d N_F1ON_MI33_g N_VDD_MI33_s ptft L=1.8e-05 W=0.00012
XMI41 N_VSS_MI41_d N_VSS_MI41_g N_net160_MI41_s ptft L=1.8e-05 W=4e-05
XMI30 N_VSS_MI41_d N_VSS_MI30_g N_net159_MI30_s ptft L=1.8e-05 W=4e-05
XMI39 N_net160_MI39_d N_F1N_MI39_g N_VDD_MI39_s ptft L=1.8e-05 W=0.00012
XMI32 N_net159_MI32_d N_F1_MI32_g N_VDD_MI32_s ptft L=1.8e-05 W=0.00012
XMI36 N_F1ON_MI36_d N_F1N_MI36_g N_VDD_MI36_s ptft L=1.8e-05 W=0.00024
XMI35 N_F1O_MI35_d N_F1_MI35_g N_VDD_MI35_s ptft L=1.8e-05 W=0.00024
XMI40 N_VSS_MI40_d N_net160_MI40_g N_F1ON_MI40_s ptft L=1.8e-05 W=0.00048
XMI31 N_VSS_MI40_d N_net159_MI31_g N_F1O_MI31_s ptft L=1.8e-05 W=0.00048
XMI37 N_F1ON_MI37_d N_F1O_MI37_g N_VDD_MI37_s ptft L=1.8e-05 W=0.00024
XMI34 N_F1O_MI34_d N_F1ON_MI34_g N_VDD_MI34_s ptft L=1.8e-05 W=0.00024
XMI59 N_net154_MI59_d N_::CK_MI59_g N_VDD_MI59_s ptft L=1.8e-05 W=0.00012
XMI53 N_net158_MI53_d N_::CK_MI53_g N_VDD_MI53_s ptft L=1.8e-05 W=0.00012
XMI56 N_VSS_MI56_d N_VSS_MI56_g N_net154_MI56_s ptft L=1.8e-05 W=4e-05
XMI50 N_VSS_MI56_d N_VSS_MI50_g N_net158_MI50_s ptft L=1.8e-05 W=4e-05
XMI58 N_net154_MI58_d N_F1ON_MI58_g N_VDD_MI58_s ptft L=1.8e-05 W=0.00012
XMI52 N_net158_MI52_d N_F1O_MI52_g N_VDD_MI52_s ptft L=1.8e-05 W=0.00012
XMI61 N_F2N_MI61_d N_F1ON_MI61_g N_VDD_MI61_s ptft L=1.8e-05 W=0.00024
XMI55 N_F2_MI55_d N_F1O_MI55_g N_VDD_MI55_s ptft L=1.8e-05 W=0.00024
XMI57 N_VSS_MI57_d N_net154_MI57_g N_F2N_MI57_s ptft L=1.8e-05 W=0.00048
XMI51 N_VSS_MI57_d N_net158_MI51_g N_F2_MI51_s ptft L=1.8e-05 W=0.00048
XMI60 N_F2N_MI60_d N_::CK_MI60_g N_VDD_MI60_s ptft L=1.8e-05 W=0.00024
XMI54 N_F2_MI54_d N_::CK_MI54_g N_VDD_MI54_s ptft L=1.8e-05 W=0.00024
XMI70 N_net153_MI70_d N_Q_MI70_g N_VDD_MI70_s ptft L=1.8e-05 W=0.00012
XMI65 N_net155_MI65_d N_QN_MI65_g N_VDD_MI65_s ptft L=1.8e-05 W=0.00012
XMI73 N_VSS_MI73_d N_VSS_MI73_g N_net153_MI73_s ptft L=1.8e-05 W=4e-05
XMI62 N_VSS_MI73_d N_VSS_MI62_g N_net155_MI62_s ptft L=1.8e-05 W=4e-05
XMI71 N_net153_MI71_d N_F2N_MI71_g N_VDD_MI71_s ptft L=1.8e-05 W=0.00012
XMI64 N_net155_MI64_d N_F2_MI64_g N_VDD_MI64_s ptft L=1.8e-05 W=0.00012
XMI68 N_QN_MI68_d N_F2N_MI68_g N_VDD_MI68_s ptft L=1.8e-05 W=0.00024
XMI67 N_Q_MI67_d N_F2_MI67_g N_VDD_MI67_s ptft L=1.8e-05 W=0.00024
XMI72 N_VSS_MI72_d N_net153_MI72_g N_QN_MI72_s ptft L=1.8e-05 W=0.00048
XMI63 N_VSS_MI72_d N_net155_MI63_g N_Q_MI63_s ptft L=1.8e-05 W=0.00048
XMI69 N_QN_MI69_d N_Q_MI69_g N_VDD_MI69_s ptft L=1.8e-05 W=0.00024
XMI66 N_Q_MI66_d N_QN_MI66_g N_VDD_MI66_s ptft L=1.8e-05 W=0.00024
*
.include "DFFD1.cdl.DFFD1.pxi"
*
.ends
*
*
