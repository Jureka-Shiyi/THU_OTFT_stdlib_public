* File: XOR2D2.cdl
* Created: Wed Jan 15 23:42:42 2025
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "/data/zhengyj/OTFT_stdlib/subckts/XOR2D2.cdl.pex"
.subckt XOR2D2  IN2 IN1 VSS VDD OUT
* 
* OUT	OUT
* VDD	VDD
* VSS	VSS
* IN1	IN1
* IN2	IN2
XMI1 N_net17_MI1_d N_IN1_MI1_g N_VSS_MI1_s ntft L=4e-06 W=4e-05
XMI15 N_net19_MI15_d N_IN2_MI15_g N_VSS_MI15_s ntft L=4e-06 W=4e-05
XMI11 N_net17_MI11_d N_net19_MI11_g N_net20_MI11_s ntft L=4e-06 W=4e-05
XMI0 N_net17_MI0_d N_IN1_MI0_g N_VDD_MI0_s ptft L=4e-06 W=2e-05
XMI14 N_net19_MI14_d N_IN2_MI14_g N_VDD_MI14_s ptft L=4e-06 W=2e-05
XMI10 N_net17_MI10_d N_IN2_MI10_g N_net20_MI10_s ptft L=4e-06 W=2e-05
XMI9 net21 N_net17_MI9_g N_VSS_MI9_s ntft L=4e-06 W=8e-05
XMI8 N_net20_MI8_d N_IN2_MI8_g net21 ntft L=4e-06 W=8e-05
XMI13 N_OUT_MI13_d N_net20_MI13_g N_VSS_MI13_s ntft L=4e-06 W=8e-05
XMI7 N_net20_MI7_d N_net19_MI7_g net18 ptft L=4e-06 W=4e-05
XMI6 net18 N_net17_MI6_g N_VDD_MI6_s ptft L=4e-06 W=4e-05
XMI12 N_OUT_MI12_d N_net20_MI12_g N_VDD_MI12_s ptft L=4e-06 W=4e-05
c_506 net21 0 0.410184f
c_518 net18 0 0.230204f
*
.include "/data/zhengyj/OTFT_stdlib/subckts/XOR2D2.cdl.XOR2D2.pxi"
*
.ends
*
*
