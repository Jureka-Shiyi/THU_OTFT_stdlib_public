* SPICE NETLIST
***************************************

.SUBCKT NAND2D8 VSS OUT VDD IN1 IN2
** N=6 EP=5 IP=0 FDC=88
M0 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=80000 $Y=430000 $D=0
M1 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=120000 $Y=430000 $D=0
M2 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=160000 $Y=430000 $D=0
M3 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=200000 $Y=430000 $D=0
M4 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=240000 $Y=430000 $D=0
M5 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=280000 $Y=430000 $D=0
M6 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=320000 $Y=430000 $D=0
M7 1 VSS VSS ptft L=1e-05 W=0.0001 $X=325400 $Y=172400 $D=0
M8 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=360000 $Y=430000 $D=0
M9 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=365400 $Y=172400 $D=0
M10 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=400000 $Y=430000 $D=0
M11 1 VSS VSS ptft L=1e-05 W=0.0001 $X=405400 $Y=172400 $D=0
M12 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=440000 $Y=430000 $D=0
M13 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=445400 $Y=172400 $D=0
M14 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=480000 $Y=430000 $D=0
M15 1 VSS VSS ptft L=1e-05 W=0.0001 $X=485400 $Y=172400 $D=0
M16 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=520000 $Y=430000 $D=0
M17 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=525400 $Y=172400 $D=0
M18 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=560000 $Y=430000 $D=0
M19 1 VSS VSS ptft L=1e-05 W=0.0001 $X=565400 $Y=172400 $D=0
M20 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=600000 $Y=430000 $D=0
M21 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=605400 $Y=172400 $D=0
M22 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=640000 $Y=430000 $D=0
M23 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=680000 $Y=430000 $D=0
M24 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=720000 $Y=43600 $D=0
M25 1 IN1 VDD ptft L=1e-05 W=0.0004 $X=720000 $Y=430000 $D=0
M26 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=760000 $Y=43600 $D=0
M27 VDD IN1 1 ptft L=1e-05 W=0.0004 $X=760000 $Y=430000 $D=0
M28 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=800000 $Y=43600 $D=0
M29 1 IN1 VDD ptft L=1e-05 W=0.0004 $X=800000 $Y=430000 $D=0
M30 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=840000 $Y=43600 $D=0
M31 VDD IN1 1 ptft L=1e-05 W=0.0004 $X=840000 $Y=430000 $D=0
M32 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=880000 $Y=43600 $D=0
M33 1 IN1 VDD ptft L=1e-05 W=0.0004 $X=880000 $Y=430000 $D=0
M34 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=920000 $Y=43600 $D=0
M35 VDD IN1 1 ptft L=1e-05 W=0.0004 $X=920000 $Y=430000 $D=0
M36 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=960000 $Y=43600 $D=0
M37 1 IN1 VDD ptft L=1e-05 W=0.0004 $X=960000 $Y=430000 $D=0
M38 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1000000 $Y=43600 $D=0
M39 VDD IN1 1 ptft L=1e-05 W=0.0004 $X=1000000 $Y=430000 $D=0
M40 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1040000 $Y=43600 $D=0
M41 1 IN2 VDD ptft L=1e-05 W=0.0004 $X=1040000 $Y=430000 $D=0
M42 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1080000 $Y=43600 $D=0
M43 VDD IN2 1 ptft L=1e-05 W=0.0004 $X=1080000 $Y=430000 $D=0
M44 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1120000 $Y=43600 $D=0
M45 1 IN2 VDD ptft L=1e-05 W=0.0004 $X=1120000 $Y=430000 $D=0
M46 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1160000 $Y=43600 $D=0
M47 VDD IN2 1 ptft L=1e-05 W=0.0004 $X=1160000 $Y=430000 $D=0
M48 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1200000 $Y=43600 $D=0
M49 1 IN2 VDD ptft L=1e-05 W=0.0004 $X=1200000 $Y=430000 $D=0
M50 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1240000 $Y=43600 $D=0
M51 VDD IN2 1 ptft L=1e-05 W=0.0004 $X=1240000 $Y=430000 $D=0
M52 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1280000 $Y=43600 $D=0
M53 1 IN2 VDD ptft L=1e-05 W=0.0004 $X=1280000 $Y=430000 $D=0
M54 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1320000 $Y=43600 $D=0
M55 VDD IN2 1 ptft L=1e-05 W=0.0004 $X=1320000 $Y=430000 $D=0
M56 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1360000 $Y=43600 $D=0
M57 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=1360000 $Y=430000 $D=0
M58 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1400000 $Y=43600 $D=0
M59 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=1400000 $Y=430000 $D=0
M60 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1440000 $Y=43600 $D=0
M61 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=1440000 $Y=430000 $D=0
M62 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1480000 $Y=43600 $D=0
M63 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=1480000 $Y=430000 $D=0
M64 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1520000 $Y=43600 $D=0
M65 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=1520000 $Y=430000 $D=0
M66 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1560000 $Y=43600 $D=0
M67 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=1560000 $Y=430000 $D=0
M68 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1600000 $Y=43600 $D=0
M69 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=1600000 $Y=430000 $D=0
M70 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1640000 $Y=43600 $D=0
M71 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=1640000 $Y=430000 $D=0
M72 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1680000 $Y=43600 $D=0
M73 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=1680000 $Y=430000 $D=0
M74 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1720000 $Y=43600 $D=0
M75 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=1720000 $Y=430000 $D=0
M76 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1760000 $Y=43600 $D=0
M77 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=1760000 $Y=430000 $D=0
M78 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1800000 $Y=43600 $D=0
M79 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=1800000 $Y=430000 $D=0
M80 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1840000 $Y=43600 $D=0
M81 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=1840000 $Y=430000 $D=0
M82 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1880000 $Y=43600 $D=0
M83 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=1880000 $Y=430000 $D=0
M84 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=1920000 $Y=43600 $D=0
M85 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=1920000 $Y=430000 $D=0
M86 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1960000 $Y=43600 $D=0
M87 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=1960000 $Y=430000 $D=0
.ENDS
***************************************
