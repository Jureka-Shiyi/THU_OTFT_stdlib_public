* File: BUFD2.cdl
* Created: Sat Dec 27 12:57:47 2025
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "BUFD2.cdl.pex"
.subckt BUFD2  VSS VDD OUT IN
* 
* IN	IN
* OUT	OUT
* VDD	VDD
* VSS	VSS
XMI5 N_VSS_MI5_d N_VSS_MI5_g N_net2_MI5_s ptft L=4e-05 W=0.0001
XMI4 N_net2_MI4_d N_IN_MI4_g N_VDD_MI4_s ptft L=1e-05 W=0.0002
XMI5@2 N_VSS_MI5@2_d N_VSS_MI5@2_g N_net2_MI5_s ptft L=4e-05 W=0.0001
XMI4@2 N_net2_MI4@2_d N_IN_MI4@2_g N_VDD_MI4_s ptft L=1e-05 W=0.0002
XMI7 N_VSS_MI7_d N_net2_MI7_g N_net1_MI7_s ptft L=1e-05 W=0.0002
XMI6 N_net1_MI6_d N_IN_MI6_g N_VDD_MI6_s ptft L=1e-05 W=0.0002
XMI7@4 N_VSS_MI7_d N_net2_MI7@4_g N_net1_MI7@4_s ptft L=1e-05 W=0.0002
XMI6@4 N_net1_MI6@4_d N_IN_MI6@4_g N_VDD_MI6_s ptft L=1e-05 W=0.0002
XMI7@3 N_VSS_MI7@3_d N_net2_MI7@3_g N_net1_MI7@4_s ptft L=1e-05 W=0.0002
XMI6@3 N_net1_MI6@4_d N_IN_MI6@3_g N_VDD_MI6@3_s ptft L=1e-05 W=0.0002
XMI7@2 N_VSS_MI7@3_d N_net2_MI7@2_g N_net1_MI7@2_s ptft L=1e-05 W=0.0002
XMI6@2 N_net1_MI6@2_d N_IN_MI6@2_g N_VDD_MI6@3_s ptft L=1e-05 W=0.0002
XMI11 N_VSS_MI11_d N_VSS_MI11_g N_net3_MI11_s ptft L=4e-05 W=0.0001
XMI9 N_net3_MI9_d N_net1_MI9_g N_VDD_MI9_s ptft L=1e-05 W=0.0002
XMI11@2 N_VSS_MI11@2_d N_VSS_MI11@2_g N_net3_MI11_s ptft L=4e-05 W=0.0001
XMI9@2 N_net3_MI9@2_d N_net1_MI9@2_g N_VDD_MI9_s ptft L=1e-05 W=0.0002
XMI10 N_VSS_MI10_d N_net3_MI10_g N_OUT_MI10_s ptft L=1e-05 W=0.0002
XMI8 N_OUT_MI8_d N_net1_MI8_g N_VDD_MI8_s ptft L=1e-05 W=0.0002
XMI10@4 N_VSS_MI10_d N_net3_MI10@4_g N_OUT_MI10@4_s ptft L=1e-05 W=0.0002
XMI8@4 N_OUT_MI8@4_d N_net1_MI8@4_g N_VDD_MI8_s ptft L=1e-05 W=0.0002
XMI10@3 N_VSS_MI10@3_d N_net3_MI10@3_g N_OUT_MI10@4_s ptft L=1e-05 W=0.0002
XMI8@3 N_OUT_MI8@4_d N_net1_MI8@3_g N_VDD_MI8@3_s ptft L=1e-05 W=0.0002
XMI10@2 N_VSS_MI10@3_d N_net3_MI10@2_g N_OUT_MI10@2_s ptft L=1e-05 W=0.0002
XMI8@2 N_OUT_MI8@2_d N_net1_MI8@2_g N_VDD_MI8@3_s ptft L=1e-05 W=0.0002
*
.include "BUFD2.cdl.BUFD2.pxi"
*
.ends
*
*
