* SPICE NETLIST
***************************************

.SUBCKT DFFD1 CK D VSS VDD QN Q
** N=26 EP=6 IP=0 FDC=60
M0 VDD 7 4 ptft L=1.8e-05 W=0.00016 $X=584500 $Y=145500 $D=0
M1 VDD CK 5 ptft L=1.8e-05 W=0.00016 $X=584500 $Y=413500 $D=0
M2 VDD D 6 ptft L=1.8e-05 W=0.00016 $X=584500 $Y=681500 $D=0
M3 4 VSS VSS ptft L=1.8e-05 W=4e-05 $X=684500 $Y=44000 $D=0
M4 5 VSS VSS ptft L=1.8e-05 W=4e-05 $X=684500 $Y=312000 $D=0
M5 6 VSS VSS ptft L=1.8e-05 W=4e-05 $X=684500 $Y=580000 $D=0
M6 18 4 VSS ptft L=1.8e-05 W=0.00032 $X=944500 $Y=85500 $D=0
M7 VDD 7 18 ptft L=1.8e-05 W=0.00032 $X=944500 $Y=145500 $D=0
M8 7 5 VSS ptft L=1.8e-05 W=0.00032 $X=944500 $Y=353500 $D=0
M9 VDD CK 7 ptft L=1.8e-05 W=0.00032 $X=944500 $Y=413500 $D=0
M10 10 6 VSS ptft L=1.8e-05 W=0.00032 $X=944500 $Y=621500 $D=0
M11 VDD D 10 ptft L=1.8e-05 W=0.00032 $X=944500 $Y=681500 $D=0
M12 8 7 VDD ptft L=1.8e-05 W=0.00012 $X=1590500 $Y=204500 $D=0
M13 VDD 7 9 ptft L=1.8e-05 W=0.00012 $X=1590500 $Y=588500 $D=0
M14 VSS VSS 8 ptft L=1.8e-05 W=4e-05 $X=1710500 $Y=362000 $D=0
M15 9 VSS VSS ptft L=1.8e-05 W=4e-05 $X=1710500 $Y=431000 $D=0
M16 8 10 VDD ptft L=1.8e-05 W=0.00012 $X=1750500 $Y=204500 $D=0
M17 VDD D 9 ptft L=1.8e-05 W=0.00012 $X=1750500 $Y=588500 $D=0
M18 15 10 VDD ptft L=1.8e-05 W=0.00024 $X=1930500 $Y=204500 $D=0
M19 VDD D 14 ptft L=1.8e-05 W=0.00024 $X=1930500 $Y=588500 $D=0
M20 VSS 8 15 ptft L=1.8e-05 W=0.00048 $X=1970500 $Y=320500 $D=0
M21 14 9 VSS ptft L=1.8e-05 W=0.00048 $X=1970500 $Y=472500 $D=0
M22 15 7 VDD ptft L=1.8e-05 W=0.00024 $X=2210500 $Y=204500 $D=0
M23 VDD 7 14 ptft L=1.8e-05 W=0.00024 $X=2210500 $Y=588500 $D=0
M24 12 17 VDD ptft L=1.8e-05 W=0.00012 $X=2556500 $Y=204500 $D=0
M25 VDD 16 13 ptft L=1.8e-05 W=0.00012 $X=2556500 $Y=588500 $D=0
M26 VSS VSS 12 ptft L=1.8e-05 W=4e-05 $X=2676500 $Y=362000 $D=0
M27 13 VSS VSS ptft L=1.8e-05 W=4e-05 $X=2676500 $Y=431000 $D=0
M28 12 15 VDD ptft L=1.8e-05 W=0.00012 $X=2716500 $Y=204500 $D=0
M29 VDD 14 13 ptft L=1.8e-05 W=0.00012 $X=2716500 $Y=588500 $D=0
M30 16 15 VDD ptft L=1.8e-05 W=0.00024 $X=2896500 $Y=204500 $D=0
M31 VDD 14 17 ptft L=1.8e-05 W=0.00024 $X=2896500 $Y=588500 $D=0
M32 VSS 12 16 ptft L=1.8e-05 W=0.00048 $X=2936500 $Y=320500 $D=0
M33 17 13 VSS ptft L=1.8e-05 W=0.00048 $X=2936500 $Y=472500 $D=0
M34 16 17 VDD ptft L=1.8e-05 W=0.00024 $X=3176500 $Y=204500 $D=0
M35 VDD 16 17 ptft L=1.8e-05 W=0.00024 $X=3176500 $Y=588500 $D=0
M36 19 18 VDD ptft L=1.8e-05 W=0.00012 $X=3690500 $Y=204500 $D=0
M37 VDD 18 20 ptft L=1.8e-05 W=0.00012 $X=3690500 $Y=588500 $D=0
M38 VSS VSS 19 ptft L=1.8e-05 W=4e-05 $X=3810500 $Y=362000 $D=0
M39 20 VSS VSS ptft L=1.8e-05 W=4e-05 $X=3810500 $Y=431000 $D=0
M40 19 16 VDD ptft L=1.8e-05 W=0.00012 $X=3850500 $Y=204500 $D=0
M41 VDD 17 20 ptft L=1.8e-05 W=0.00012 $X=3850500 $Y=588500 $D=0
M42 23 16 VDD ptft L=1.8e-05 W=0.00024 $X=4030500 $Y=204500 $D=0
M43 VDD 17 24 ptft L=1.8e-05 W=0.00024 $X=4030500 $Y=588500 $D=0
M44 VSS 19 23 ptft L=1.8e-05 W=0.00048 $X=4070500 $Y=320500 $D=0
M45 24 20 VSS ptft L=1.8e-05 W=0.00048 $X=4070500 $Y=472500 $D=0
M46 23 18 VDD ptft L=1.8e-05 W=0.00024 $X=4310500 $Y=204500 $D=0
M47 VDD 18 24 ptft L=1.8e-05 W=0.00024 $X=4310500 $Y=588500 $D=0
M48 21 Q VDD ptft L=1.8e-05 W=0.00012 $X=4656500 $Y=204500 $D=0
M49 VDD QN 22 ptft L=1.8e-05 W=0.00012 $X=4656500 $Y=588500 $D=0
M50 VSS VSS 21 ptft L=1.8e-05 W=4e-05 $X=4776500 $Y=362000 $D=0
M51 22 VSS VSS ptft L=1.8e-05 W=4e-05 $X=4776500 $Y=431000 $D=0
M52 21 23 VDD ptft L=1.8e-05 W=0.00012 $X=4816500 $Y=204500 $D=0
M53 VDD 24 22 ptft L=1.8e-05 W=0.00012 $X=4816500 $Y=588500 $D=0
M54 QN 23 VDD ptft L=1.8e-05 W=0.00024 $X=4996500 $Y=204500 $D=0
M55 VDD 24 Q ptft L=1.8e-05 W=0.00024 $X=4996500 $Y=588500 $D=0
M56 VSS 21 QN ptft L=1.8e-05 W=0.00048 $X=5036500 $Y=320500 $D=0
M57 Q 22 VSS ptft L=1.8e-05 W=0.00048 $X=5036500 $Y=472500 $D=0
M58 QN Q VDD ptft L=1.8e-05 W=0.00024 $X=5276500 $Y=204500 $D=0
M59 VDD QN Q ptft L=1.8e-05 W=0.00024 $X=5276500 $Y=588500 $D=0
.ENDS
***************************************
