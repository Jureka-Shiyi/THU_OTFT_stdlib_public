* SPICE NETLIST
***************************************

.SUBCKT BUFD2 VSS VDD OUT IN
** N=7 EP=4 IP=0 FDC=24
M0 1 VSS VSS ptft L=4e-05 W=0.0001 $X=112000 $Y=300000 $D=0
M1 VDD IN 1 ptft L=1e-05 W=0.0002 $X=142000 $Y=580000 $D=0
M2 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=192000 $Y=300000 $D=0
M3 1 IN VDD ptft L=1e-05 W=0.0002 $X=192000 $Y=580000 $D=0
M4 VSS 1 3 ptft L=1e-05 W=0.0002 $X=362000 $Y=180000 $D=0
M5 VDD IN 3 ptft L=1e-05 W=0.0002 $X=362000 $Y=580000 $D=0
M6 3 1 VSS ptft L=1e-05 W=0.0002 $X=412000 $Y=180000 $D=0
M7 3 IN VDD ptft L=1e-05 W=0.0002 $X=412000 $Y=580000 $D=0
M8 VSS 1 3 ptft L=1e-05 W=0.0002 $X=462000 $Y=180000 $D=0
M9 VDD IN 3 ptft L=1e-05 W=0.0002 $X=462000 $Y=580000 $D=0
M10 3 1 VSS ptft L=1e-05 W=0.0002 $X=512000 $Y=180000 $D=0
M11 3 IN VDD ptft L=1e-05 W=0.0002 $X=512000 $Y=580000 $D=0
M12 4 VSS VSS ptft L=4e-05 W=0.0001 $X=704000 $Y=300000 $D=0
M13 VDD 3 4 ptft L=1e-05 W=0.0002 $X=734000 $Y=580000 $D=0
M14 VSS VSS 4 ptft L=4e-05 W=0.0001 $X=784000 $Y=300000 $D=0
M15 4 3 VDD ptft L=1e-05 W=0.0002 $X=784000 $Y=580000 $D=0
M16 VSS 4 OUT ptft L=1e-05 W=0.0002 $X=954000 $Y=180000 $D=0
M17 VDD 3 OUT ptft L=1e-05 W=0.0002 $X=954000 $Y=580000 $D=0
M18 OUT 4 VSS ptft L=1e-05 W=0.0002 $X=1004000 $Y=180000 $D=0
M19 OUT 3 VDD ptft L=1e-05 W=0.0002 $X=1004000 $Y=580000 $D=0
M20 VSS 4 OUT ptft L=1e-05 W=0.0002 $X=1054000 $Y=180000 $D=0
M21 VDD 3 OUT ptft L=1e-05 W=0.0002 $X=1054000 $Y=580000 $D=0
M22 OUT 4 VSS ptft L=1e-05 W=0.0002 $X=1104000 $Y=180000 $D=0
M23 OUT 3 VDD ptft L=1e-05 W=0.0002 $X=1104000 $Y=580000 $D=0
.ENDS
***************************************
