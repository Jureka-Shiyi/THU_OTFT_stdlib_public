* SPICE NETLIST
***************************************

.SUBCKT INVD4 VSS VDD OUT IN
** N=5 EP=4 IP=0 FDC=24
M0 1 VSS VSS ptft L=4e-05 W=0.0001 $X=68000 $Y=300000 $D=0
M1 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=148000 $Y=300000 $D=0
M2 VDD IN 1 ptft L=1e-05 W=0.0002 $X=158000 $Y=580000 $D=0
M3 1 IN VDD ptft L=1e-05 W=0.0002 $X=208000 $Y=580000 $D=0
M4 1 VSS VSS ptft L=4e-05 W=0.0001 $X=228000 $Y=300000 $D=0
M5 VDD IN 1 ptft L=1e-05 W=0.0002 $X=258000 $Y=580000 $D=0
M6 VSS VSS 1 ptft L=4e-05 W=0.0001 $X=308000 $Y=300000 $D=0
M7 1 IN VDD ptft L=1e-05 W=0.0002 $X=308000 $Y=580000 $D=0
M8 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=478000 $Y=180000 $D=0
M9 VDD IN OUT ptft L=1e-05 W=0.0002 $X=478000 $Y=580000 $D=0
M10 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=528000 $Y=180000 $D=0
M11 OUT IN VDD ptft L=1e-05 W=0.0002 $X=528000 $Y=580000 $D=0
M12 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=578000 $Y=180000 $D=0
M13 VDD IN OUT ptft L=1e-05 W=0.0002 $X=578000 $Y=580000 $D=0
M14 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=628000 $Y=180000 $D=0
M15 OUT IN VDD ptft L=1e-05 W=0.0002 $X=628000 $Y=580000 $D=0
M16 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=678000 $Y=180000 $D=0
M17 VDD IN OUT ptft L=1e-05 W=0.0002 $X=678000 $Y=580000 $D=0
M18 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=728000 $Y=180000 $D=0
M19 OUT IN VDD ptft L=1e-05 W=0.0002 $X=728000 $Y=580000 $D=0
M20 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=778000 $Y=180000 $D=0
M21 VDD IN OUT ptft L=1e-05 W=0.0002 $X=778000 $Y=580000 $D=0
M22 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=828000 $Y=180000 $D=0
M23 OUT IN VDD ptft L=1e-05 W=0.0002 $X=828000 $Y=580000 $D=0
.ENDS
***************************************
