* SPICE NETLIST
***************************************

.SUBCKT NAND2D4 VSS OUT VDD IN1 IN2
** N=6 EP=5 IP=0 FDC=44
M0 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=80000 $Y=430000 $D=0
M1 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=120000 $Y=430000 $D=0
M2 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=160000 $Y=430000 $D=0
M3 1 VSS VSS ptft L=1e-05 W=0.0001 $X=165400 $Y=172400 $D=0
M4 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=200000 $Y=430000 $D=0
M5 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=205400 $Y=172400 $D=0
M6 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=240000 $Y=430000 $D=0
M7 1 VSS VSS ptft L=1e-05 W=0.0001 $X=245400 $Y=172400 $D=0
M8 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=280000 $Y=430000 $D=0
M9 VSS VSS 1 ptft L=1e-05 W=0.0001 $X=285400 $Y=172400 $D=0
M10 OUT IN1 VDD ptft L=1e-05 W=0.0004 $X=320000 $Y=430000 $D=0
M11 VDD IN1 OUT ptft L=1e-05 W=0.0004 $X=360000 $Y=430000 $D=0
M12 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=400000 $Y=43600 $D=0
M13 1 IN1 VDD ptft L=1e-05 W=0.0004 $X=400000 $Y=430000 $D=0
M14 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=440000 $Y=43600 $D=0
M15 VDD IN1 1 ptft L=1e-05 W=0.0004 $X=440000 $Y=430000 $D=0
M16 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=480000 $Y=43600 $D=0
M17 1 IN1 VDD ptft L=1e-05 W=0.0004 $X=480000 $Y=430000 $D=0
M18 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=520000 $Y=43600 $D=0
M19 VDD IN1 1 ptft L=1e-05 W=0.0004 $X=520000 $Y=430000 $D=0
M20 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=560000 $Y=43600 $D=0
M21 1 IN2 VDD ptft L=1e-05 W=0.0004 $X=560000 $Y=430000 $D=0
M22 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=600000 $Y=43600 $D=0
M23 VDD IN2 1 ptft L=1e-05 W=0.0004 $X=600000 $Y=430000 $D=0
M24 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=640000 $Y=43600 $D=0
M25 1 IN2 VDD ptft L=1e-05 W=0.0004 $X=640000 $Y=430000 $D=0
M26 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=680000 $Y=43600 $D=0
M27 VDD IN2 1 ptft L=1e-05 W=0.0004 $X=680000 $Y=430000 $D=0
M28 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=720000 $Y=43600 $D=0
M29 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=720000 $Y=430000 $D=0
M30 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=760000 $Y=43600 $D=0
M31 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=760000 $Y=430000 $D=0
M32 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=800000 $Y=43600 $D=0
M33 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=800000 $Y=430000 $D=0
M34 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=840000 $Y=43600 $D=0
M35 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=840000 $Y=430000 $D=0
M36 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=880000 $Y=43600 $D=0
M37 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=880000 $Y=430000 $D=0
M38 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=920000 $Y=43600 $D=0
M39 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=920000 $Y=430000 $D=0
M40 OUT 1 VSS ptft L=1e-05 W=0.0002 $X=960000 $Y=43600 $D=0
M41 OUT IN2 VDD ptft L=1e-05 W=0.0004 $X=960000 $Y=430000 $D=0
M42 VSS 1 OUT ptft L=1e-05 W=0.0002 $X=1000000 $Y=43600 $D=0
M43 VDD IN2 OUT ptft L=1e-05 W=0.0004 $X=1000000 $Y=430000 $D=0
.ENDS
***************************************
