* File: INVD16.cdl
* Created: Sat Aug 17 14:52:21 2024
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "/data/zhengyj/OTFT_stdlib/subckts/INVD16.cdl.pex"
.subckt INVD16  IN OUT VDD VSS
* 
* VSS	VSS
* VDD	VDD
* OUT	OUT
* IN	IN
XMI6 N_OUT_MI6_d N_IN_MI6_g N_VDD_MI6_s ptft L=4e-06 W=8e-05
XMI6@2 N_OUT_MI6_d N_IN_MI6@2_g N_VDD_MI6@2_s ptft L=4e-06 W=8e-05
XMI0 N_OUT_MI0_d N_IN_MI0_g N_VSS_MI0_s ntft L=4e-06 W=8e-05
XMI1@2 N_OUT_MI0_d N_IN_MI1@2_g N_VSS_MI1@2_s ntft L=4e-06 W=8e-05
XMI1 N_OUT_MI1_d N_IN_MI1_g N_VSS_MI1_s ntft L=4e-06 W=8e-05
XMI0@2 N_OUT_MI1_d N_IN_MI0@2_g N_VSS_MI0@2_s ntft L=4e-06 W=8e-05
*
.include "/data/zhengyj/OTFT_stdlib/subckts/INVD16.cdl.INVD16.pxi"
*
.ends
*
*
