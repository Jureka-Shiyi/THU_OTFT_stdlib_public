* SPICE NETLIST
***************************************

.SUBCKT NOR2D1 VSS VDD OUT IN2 IN1
** N=8 EP=5 IP=0 FDC=18
M0 1 VSS VSS ptft L=1e-05 W=0.0001 $X=90000 $Y=160000 $D=0
M1 1 IN2 3 ptft L=1e-05 W=0.0002 $X=100000 $Y=310000 $D=0
M2 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=100000 $Y=630000 $D=0
M3 3 IN2 1 ptft L=1e-05 W=0.0002 $X=140000 $Y=310000 $D=0
M4 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=140000 $Y=630000 $D=0
M5 1 IN2 3 ptft L=1e-05 W=0.0002 $X=180000 $Y=310000 $D=0
M6 VDD IN1 3 ptft L=1e-05 W=0.0002 $X=180000 $Y=630000 $D=0
M7 3 IN2 1 ptft L=1e-05 W=0.0002 $X=220000 $Y=310000 $D=0
M8 3 IN1 VDD ptft L=1e-05 W=0.0002 $X=220000 $Y=630000 $D=0
M9 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=330000 $Y=310000 $D=0
M10 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=330000 $Y=630000 $D=0
M11 OUT 1 VSS ptft L=1e-05 W=0.0001 $X=355000 $Y=120000 $D=0
M12 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=370000 $Y=310000 $D=0
M13 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=370000 $Y=630000 $D=0
M14 OUT IN2 6 ptft L=1e-05 W=0.0002 $X=410000 $Y=310000 $D=0
M15 VDD IN1 6 ptft L=1e-05 W=0.0002 $X=410000 $Y=630000 $D=0
M16 6 IN2 OUT ptft L=1e-05 W=0.0002 $X=450000 $Y=310000 $D=0
M17 6 IN1 VDD ptft L=1e-05 W=0.0002 $X=450000 $Y=630000 $D=0
.ENDS
***************************************
