* File: AND2D8.cdl
* Created: Wed Jan 15 18:48:53 2025
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "/data/zhengyj/OTFT_stdlib/subckts/AND2D8.cdl.pex"
.subckt AND2D8  IN1 IN2 VDD VSS OUT
* 
* OUT	OUT
* VSS	VSS
* VDD	VDD
* IN2	IN2
* IN1	IN1
XMI0 N_net11_MI0_d N_IN1_MI0_g N_VDD_MI0_s ptft L=4e-06 W=8e-05
XMI1 N_net11_MI1_d N_IN2_MI1_g N_VDD_MI1_s ptft L=4e-06 W=8e-05
XMI9 N_OUT_MI9_d N_net11_MI9_g N_VDD_MI9_s ptft L=4e-06 W=8e-05
XMI4 N_OUT_MI4_d N_net11_MI4_g N_VDD_MI4_s ptft L=4e-06 W=8e-05
XMI3 N_net12_MI3_d N_IN1_MI3_g N_VSS_MI3_s ntft L=4e-06 W=8e-05
XMI6@2 N_net12_MI3_d N_IN1_MI6@2_g N_VSS_MI6@2_s ntft L=4e-06 W=8e-05
XMI6 N_net12_MI6_d N_IN1_MI6_g N_VSS_MI6_s ntft L=4e-06 W=8e-05
XMI3@2 N_net12_MI6_d N_IN1_MI3@2_g N_VSS_MI3@2_s ntft L=4e-06 W=8e-05
XMI8 N_net11_MI8_d N_IN2_MI8_g N_net12_MI8_s ntft L=4e-06 W=8e-05
XMI7@2 N_net11_MI7@2_d N_IN2_MI7@2_g N_net12_MI8_s ntft L=4e-06 W=8e-05
XMI7 N_net11_MI7_d N_IN2_MI7_g N_net12_MI7_s ntft L=4e-06 W=8e-05
XMI8@2 N_net11_MI8@2_d N_IN2_MI8@2_g N_net12_MI7_s ntft L=4e-06 W=8e-05
XMI2 N_OUT_MI2_d N_net11_MI2_g N_VSS_MI2_s ntft L=4e-06 W=8e-05
XMI5@2 N_OUT_MI2_d N_net11_MI5@2_g N_VSS_MI5@2_s ntft L=4e-06 W=8e-05
XMI5 N_OUT_MI5_d N_net11_MI5_g N_VSS_MI5_s ntft L=4e-06 W=8e-05
XMI2@2 N_OUT_MI5_d N_net11_MI2@2_g N_VSS_MI2@2_s ntft L=4e-06 W=8e-05
*
.include "/data/zhengyj/OTFT_stdlib/subckts/AND2D8.cdl.AND2D8.pxi"
*
.ends
*
*
