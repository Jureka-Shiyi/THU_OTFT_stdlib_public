* File: NAND2D4.cdl
* Created: Mon Dec 22 20:55:38 2025
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "NAND2D4.cdl.pex"
.subckt NAND2D4  VSS OUT VDD IN1 IN2
* 
* IN2	IN2
* IN1	IN1
* VDD	VDD
* OUT	OUT
* VSS	VSS
XMI4 N_OUT_MI4_d N_IN1_MI4_g N_VDD_MI4_s ptft L=1e-05 W=0.0004
XMI4@8 N_OUT_MI4_d N_IN1_MI4@8_g N_VDD_MI4@8_s ptft L=1e-05 W=0.0004
XMI4@7 N_OUT_MI4@7_d N_IN1_MI4@7_g N_VDD_MI4@8_s ptft L=1e-05 W=0.0004
XMI2 N_VSS_MI2_d N_VSS_MI2_g N_net14_MI2_s ptft L=1e-05 W=0.0001
XMI4@6 N_OUT_MI4@7_d N_IN1_MI4@6_g N_VDD_MI4@6_s ptft L=1e-05 W=0.0004
XMI2@4 N_VSS_MI2@4_d N_VSS_MI2@4_g N_net14_MI2_s ptft L=1e-05 W=0.0001
XMI4@5 N_OUT_MI4@5_d N_IN1_MI4@5_g N_VDD_MI4@6_s ptft L=1e-05 W=0.0004
XMI2@3 N_VSS_MI2@4_d N_VSS_MI2@3_g N_net14_MI2@3_s ptft L=1e-05 W=0.0001
XMI4@4 N_OUT_MI4@5_d N_IN1_MI4@4_g N_VDD_MI4@4_s ptft L=1e-05 W=0.0004
XMI2@2 N_VSS_MI2@2_d N_VSS_MI2@2_g N_net14_MI2@3_s ptft L=1e-05 W=0.0001
XMI4@3 N_OUT_MI4@3_d N_IN1_MI4@3_g N_VDD_MI4@4_s ptft L=1e-05 W=0.0004
XMI4@2 N_OUT_MI4@3_d N_IN1_MI4@2_g N_VDD_MI4@2_s ptft L=1e-05 W=0.0004
XMI5 N_VSS_MI5_d N_net14_MI5_g N_OUT_MI5_s ptft L=1e-05 W=0.0002
XMI0 N_net14_MI0_d N_IN1_MI0_g N_VDD_MI4@2_s ptft L=1e-05 W=0.0004
XMI5@16 N_VSS_MI5@16_d N_net14_MI5@16_g N_OUT_MI5_s ptft L=1e-05 W=0.0002
XMI0@4 N_net14_MI0_d N_IN1_MI0@4_g N_VDD_MI0@4_s ptft L=1e-05 W=0.0004
XMI5@15 N_VSS_MI5@16_d N_net14_MI5@15_g N_OUT_MI5@15_s ptft L=1e-05 W=0.0002
XMI0@3 N_net14_MI0@3_d N_IN1_MI0@3_g N_VDD_MI0@4_s ptft L=1e-05 W=0.0004
XMI5@14 N_VSS_MI5@14_d N_net14_MI5@14_g N_OUT_MI5@15_s ptft L=1e-05 W=0.0002
XMI0@2 N_net14_MI0@3_d N_IN1_MI0@2_g N_VDD_MI0@2_s ptft L=1e-05 W=0.0004
XMI5@13 N_VSS_MI5@14_d N_net14_MI5@13_g N_OUT_MI5@13_s ptft L=1e-05 W=0.0002
XMI1 N_net14_MI1_d N_IN2_MI1_g N_VDD_MI0@2_s ptft L=1e-05 W=0.0004
XMI5@12 N_VSS_MI5@12_d N_net14_MI5@12_g N_OUT_MI5@13_s ptft L=1e-05 W=0.0002
XMI1@4 N_net14_MI1_d N_IN2_MI1@4_g N_VDD_MI1@4_s ptft L=1e-05 W=0.0004
XMI5@11 N_VSS_MI5@12_d N_net14_MI5@11_g N_OUT_MI5@11_s ptft L=1e-05 W=0.0002
XMI1@3 N_net14_MI1@3_d N_IN2_MI1@3_g N_VDD_MI1@4_s ptft L=1e-05 W=0.0004
XMI5@10 N_VSS_MI5@10_d N_net14_MI5@10_g N_OUT_MI5@11_s ptft L=1e-05 W=0.0002
XMI1@2 N_net14_MI1@3_d N_IN2_MI1@2_g N_VDD_MI1@2_s ptft L=1e-05 W=0.0004
XMI5@9 N_VSS_MI5@10_d N_net14_MI5@9_g N_OUT_MI5@9_s ptft L=1e-05 W=0.0002
XMI3 N_OUT_MI3_d N_IN2_MI3_g N_VDD_MI1@2_s ptft L=1e-05 W=0.0004
XMI5@8 N_VSS_MI5@8_d N_net14_MI5@8_g N_OUT_MI5@9_s ptft L=1e-05 W=0.0002
XMI3@8 N_OUT_MI3_d N_IN2_MI3@8_g N_VDD_MI3@8_s ptft L=1e-05 W=0.0004
XMI5@7 N_VSS_MI5@8_d N_net14_MI5@7_g N_OUT_MI5@7_s ptft L=1e-05 W=0.0002
XMI3@7 N_OUT_MI3@7_d N_IN2_MI3@7_g N_VDD_MI3@8_s ptft L=1e-05 W=0.0004
XMI5@6 N_VSS_MI5@6_d N_net14_MI5@6_g N_OUT_MI5@7_s ptft L=1e-05 W=0.0002
XMI3@6 N_OUT_MI3@7_d N_IN2_MI3@6_g N_VDD_MI3@6_s ptft L=1e-05 W=0.0004
XMI5@5 N_VSS_MI5@6_d N_net14_MI5@5_g N_OUT_MI5@5_s ptft L=1e-05 W=0.0002
XMI3@5 N_OUT_MI3@5_d N_IN2_MI3@5_g N_VDD_MI3@6_s ptft L=1e-05 W=0.0004
XMI5@4 N_VSS_MI5@4_d N_net14_MI5@4_g N_OUT_MI5@5_s ptft L=1e-05 W=0.0002
XMI3@4 N_OUT_MI3@5_d N_IN2_MI3@4_g N_VDD_MI3@4_s ptft L=1e-05 W=0.0004
XMI5@3 N_VSS_MI5@4_d N_net14_MI5@3_g N_OUT_MI5@3_s ptft L=1e-05 W=0.0002
XMI3@3 N_OUT_MI3@3_d N_IN2_MI3@3_g N_VDD_MI3@4_s ptft L=1e-05 W=0.0004
XMI5@2 N_VSS_MI5@2_d N_net14_MI5@2_g N_OUT_MI5@3_s ptft L=1e-05 W=0.0002
XMI3@2 N_OUT_MI3@3_d N_IN2_MI3@2_g N_VDD_MI3@2_s ptft L=1e-05 W=0.0004
*
.include "NAND2D4.cdl.NAND2D4.pxi"
*
.ends
*
*
