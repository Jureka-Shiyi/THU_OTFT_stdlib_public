* File: BUFD8.cdl
* Created: Fri Dec  6 22:29:38 2024
* Program "Calibre xRC"
* Version "v2023.1_18.8"
* 
.include "/data/zhengyj/OTFT_stdlib/subckts/BUFD8.cdl.pex"
.subckt BUFD8  IN VDD OUT VSS
* 
* VSS	VSS
* OUT	OUT
* VDD	VDD
* IN	IN
XMI1 N_net1_MI1_d N_IN_MI1_g N_VSS_MI1_s ntft L=4e-06 W=8e-05
XMI0 N_net1_MI0_d N_IN_MI0_g N_VDD_MI0_s ptft L=4e-06 W=4e-05
XMI2 N_OUT_MI2_d N_net1_MI2_g N_VDD_MI2_s ptft L=4e-06 W=6e-05
XMI2@2 N_OUT_MI2_d N_net1_MI2@2_g N_VDD_MI2@2_s ptft L=4e-06 W=6e-05
XMI4 N_OUT_MI4_d N_net1_MI4_g N_VSS_MI4_s ntft L=4e-06 W=6e-05
XMI3@2 N_OUT_MI4_d N_net1_MI3@2_g N_VSS_MI3@2_s ntft L=4e-06 W=6e-05
XMI3 N_OUT_MI3_d N_net1_MI3_g N_VSS_MI3_s ntft L=4e-06 W=6e-05
XMI4@2 N_OUT_MI3_d N_net1_MI4@2_g N_VSS_MI4@2_s ntft L=4e-06 W=6e-05
*
.include "/data/zhengyj/OTFT_stdlib/subckts/BUFD8.cdl.BUFD8.pxi"
*
.ends
*
*
