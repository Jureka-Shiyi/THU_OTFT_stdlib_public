VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BOUNDARY_LEFT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BOUNDARY_LEFT 0 0 ;
  SIZE 10 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 870 10 900 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 10 30 ;
    END
  END VSS
END BOUNDARY_LEFT

MACRO BOUNDARY_RIGHT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BOUNDARY_RIGHT 0 0 ;
  SIZE 10 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 870 10 900 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 10 30 ;
    END
  END VSS
END BOUNDARY_RIGHT

MACRO DFFD1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFD1 0 0 ;
  SIZE 5700 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57 698.5 242 736.5 ;
      LAYER M1 ;
        RECT 0 702 152 732 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 30 430.5 242 468.5 ;
      LAYER M1 ;
        RECT 0 434 141.5 464 ;
    END
  END CK
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 2326 170 2591.5 210 ;
        RECT 2326 654 2613 694 ;
        RECT 3278.5 170 3562 210 ;
        RECT 4422.5 654 4701 694 ;
        RECT 4413.5 170 4702.5 210 ;
      LAYER M1 ;
        POLYGON 3382 220 3372 220 3372 231 3132 231 3132 220 3092 220 3092 231 2852 231 2852 220 2792 220 2792 231 2672 231 2672 220 2632 220 2632 231 2512 231 2512 220 2502 220 2502 170 2591.5 170 2591.5 190 3282.5 190 3282.5 170 3382 170 ;
        POLYGON 4516 694 4422.5 694 4422.5 674 2607.5 674 2607.5 694 2502 694 2502 644 2512 644 2512 633 2632 633 2632 644 2672 644 2672 633 2792 633 2792 644 2852 644 2852 633 3092 633 3092 644 3132 644 3132 633 3372 633 3372 644 3646 644 3646 633 3766 633 3766 644 3806 644 3806 633 3926 633 3926 644 3986 644 3986 633 4226 633 4226 644 4266 644 4266 633 4506 633 4506 644 4516 644 ;
        POLYGON 4516 220 4506 220 4506 231 4266 231 4266 220 4226 220 4226 231 3986 231 3986 220 3926 220 3926 231 3806 231 3806 220 3766 220 3766 231 3646 231 3646 220 3458 220 3458 170 3557.5 170 3557.5 190 4409.5 190 4409.5 170 4516 170 ;
        POLYGON 5472 231 5232 231 5232 220 5192 220 5192 231 4952 231 4952 220 4892 220 4892 231 4772 231 4772 220 4732 220 4732 231 4612 231 4612 220 4602 220 4602 170 4706 170 4706 190 5472 190 ;
        POLYGON 5482 674 4698.5 674 4698.5 694 4602 694 4602 644 4612 644 4612 633 4732 633 4732 644 4772 644 4772 633 4892 633 4892 644 4952 644 4952 633 5192 633 5192 644 5232 644 5232 633 5472 633 5472 644 5482 644 ;
        POLYGON 5700 900 0 900 0 870 182 870 182 752 311 752 311 216 540 216 540 190 700 190 700 216 900 216 900 190 1220 190 1220 216 1230 216 1230 246 341 246 341 484 540 484 540 458 700 458 700 484 900 484 900 458 1220 458 1220 484 1230 484 1230 514 341 514 341 752 540 752 540 726 700 726 700 752 900 752 900 726 1220 726 1220 752 1506 752 1506 674 1391 674 1391 190 2326 190 2326 170 2416 170 2416 220 2406 220 2406 231 2166 231 2166 220 2126 220 2126 231 1886 231 1886 220 1826 220 1826 231 1706 231 1706 220 1666 220 1666 231 1546 231 1546 220 1421 220 1421 644 1546 644 1546 633 1666 633 1666 644 1706 644 1706 633 1826 633 1826 644 1886 644 1886 633 2126 633 2126 644 2166 644 2166 633 2406 633 2406 644 2416 644 2416 694 2326 694 2326 674 1536 674 1536 782 225 782 225 870 5700 870 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 1482 555 637 555 637 634 540 634 540 596 282 596 282 822 374 822 374 852 252 852 252 30 637 30 637 98 540 98 540 60 282 60 282 298 637 298 637 366 540 366 540 328 282 328 282 566 540 566 540 525 1452 525 1452 409 1482 409 ;
        RECT 1566 379 1663 485 ;
        RECT 2532 379 2629 485 ;
        POLYGON 3643 732 3518 732 3518 414.5 3569.5 414.5 3569.5 692 3643 692 ;
        RECT 3666 379 3763 485 ;
        RECT 4632 379 4729 485 ;
      LAYER M1 ;
        POLYGON 1230 596 1220 596 1220 648 900 648 900 596 680 596 680 606.5 640 606.5 640 596 510 596 510 566 1230 566 ;
        POLYGON 1230 328 1220 328 1220 380 900 380 900 328 680 328 680 338.5 640 338.5 640 328 510 328 510 298 1230 298 ;
        POLYGON 3382 447 3372 447 3372 499 2892 499 2892 447 2672 447 2672 457.5 2632 457.5 2632 447 2406 447 2406 499 1926 499 1926 447 1706 447 1706 457.5 1666 457.5 1666 447 1482 447 1482 512 1452 512 1452 417 1666 417 1666 406.5 1706 406.5 1706 417 1926 417 1926 365 2406 365 2406 417 2632 417 2632 406.5 2672 406.5 2672 417 2892 417 2892 365 3372 365 3372 417 3382 417 ;
        POLYGON 3636 732 3442 732 3442 852 248.5 852 248.5 822 3412 822 3412 699.5 3636 699.5 ;
        POLYGON 5482 447 5472 447 5472 499 4992 499 4992 447 4772 447 4772 457.5 4732 457.5 4732 447 4506 447 4506 499 4026 499 4026 447 3806 447 3806 457.5 3766 457.5 3766 447 3570.5 447 3570.5 485 3516.5 485 3516.5 412 3570.5 412 3570.5 417 3766 417 3766 406.5 3806 406.5 3806 417 4026 417 4026 365 4506 365 4506 417 4732 417 4732 406.5 4772 406.5 4772 417 4992 417 4992 365 5472 365 5472 417 5482 417 ;
        POLYGON 5700 30 1230 30 1230 60 1220 60 1220 112 900 112 900 60 680 60 680 70.5 640 70.5 640 60 510 60 510 30 0 30 0 0 5700 0 ;
    END
  END VSS
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        POLYGON 5671 351.5 5633 351.5 5633 314 5549.5 314 5549.5 276.5 5671 276.5 ;
      LAYER M1 ;
        POLYGON 5667 547 5462 547 5462 603 5472 603 5472 615 5232 615 5232 609 5192 609 5192 615 4952 615 4952 579 5322 579 5322 529 4992 529 4992 517 5637 517 5637 280 5667 280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5498 347 5535.5 517 ;
      LAYER M1 ;
        POLYGON 5532 428.5 5502 428.5 5502 347 4992 347 4992 335 5322 335 5322 285 4952 285 4952 249 5192 249 5192 255 5232 255 5232 249 5472 249 5472 261 5462 261 5462 317 5502 317 5502 175.5 5532 175.5 ;
    END
  END QN
  OBS
    LAYER M1 ;
      POLYGON 4982.5 142 4572 142 4572 279 4496 279 4496 335 4506 335 4506 347 4026 347 4026 335 4356 335 4356 285 3986 285 3986 249 4226 249 4226 255 4266 255 4266 249 4542 249 4542 112 4982.5 112 ;
      POLYGON 4981 752 4542 752 4542 615 4266 615 4266 609 4226 609 4226 615 3986 615 3986 579 4356 579 4356 529 4026 529 4026 517 4506 517 4506 529 4496 529 4496 585 4572 585 4572 722 4981 722 ;
      POLYGON 4892 285 4662 285 4662 325.5 4772 325.5 4772 388.5 4732 388.5 4732 360 4632 360 4632 285 4612 285 4612 249 4732 249 4732 255 4772 255 4772 249 4892 249 ;
      POLYGON 4892 615 4772 615 4772 609 4732 609 4732 615 4612 615 4612 579 4632 579 4632 504 4732 504 4732 475.5 4772 475.5 4772 538.5 4662 538.5 4662 579 4892 579 ;
      POLYGON 3926 285 3696 285 3696 325.5 3806 325.5 3806 388.5 3766 388.5 3766 360 3666 360 3666 285 3646 285 3646 249 3766 249 3766 255 3806 255 3806 249 3926 249 ;
      POLYGON 3926 615 3806 615 3806 609 3766 609 3766 615 3646 615 3646 579 3666 579 3666 504 3766 504 3766 475.5 3806 475.5 3806 538.5 3696 538.5 3696 579 3926 579 ;
      POLYGON 3912 142 3432 142 3432 424.5 3402 424.5 3402 347 2892 347 2892 335 3222 335 3222 285 2852 285 2852 249 3092 249 3092 255 3132 255 3132 249 3372 249 3372 261 3362 261 3362 317 3402 317 3402 112 3912 112 ;
      POLYGON 3729.5 99.5 1288 99.5 1288 160 1220 160 1220 172 900 172 900 130 1258 130 1258 61.5 3729.5 61.5 ;
      POLYGON 3492 623.5 3462 623.5 3462 547 3362 547 3362 603 3372 603 3372 615 3132 615 3132 609 3092 609 3092 615 2852 615 2852 579 3222 579 3222 529 2892 529 2892 517 3462 517 3462 317 3492 317 ;
      POLYGON 2876.5 142 2472 142 2472 279 2396 279 2396 335 2406 335 2406 347 1926 347 1926 335 2256 335 2256 285 1886 285 1886 249 2126 249 2126 255 2166 255 2166 249 2442 249 2442 112 2876.5 112 ;
      POLYGON 2862 752 2442 752 2442 615 2166 615 2166 609 2126 609 2126 615 1886 615 1886 579 2256 579 2256 529 1926 529 1926 517 2406 517 2406 529 2396 529 2396 585 2472 585 2472 722 2862 722 ;
      POLYGON 2792 285 2562 285 2562 325.5 2672 325.5 2672 388.5 2632 388.5 2632 360 2532 360 2532 285 2512 285 2512 249 2632 249 2632 255 2672 255 2672 249 2792 249 ;
      POLYGON 2792 615 2672 615 2672 609 2632 609 2632 615 2512 615 2512 579 2532 579 2532 504 2632 504 2632 475.5 2672 475.5 2672 538.5 2562 538.5 2562 579 2792 579 ;
      POLYGON 1826 285 1596 285 1596 325.5 1706 325.5 1706 388.5 1666 388.5 1666 360 1566 360 1566 285 1546 285 1546 249 1666 249 1666 255 1706 255 1706 249 1826 249 ;
      POLYGON 1826 615 1706 615 1706 609 1666 609 1666 615 1546 615 1546 579 1566 579 1566 504 1666 504 1666 475.5 1706 475.5 1706 538.5 1596 538.5 1596 579 1826 579 ;
      POLYGON 1811.5 152.5 1343 152.5 1343 696 1220 696 1220 708 900 708 900 666 1313 666 1313 122.5 1811.5 122.5 ;
      POLYGON 1292 467 1262 467 1262 428 1220 428 1220 440 900 440 900 398 1262 398 1262 369.5 1292 369.5 ;
      POLYGON 700 172 540 172 540 117 640 117 640 88.5 680 88.5 680 160 700 160 ;
      POLYGON 700 440 540 440 540 385 640 385 640 356.5 680 356.5 680 428 700 428 ;
      POLYGON 700 708 540 708 540 653 640 653 640 624.5 680 624.5 680 696 700 696 ;
    LAYER Via1 ;
      RECT 5644.5 289 5659.5 304 ;
      RECT 5644.5 309 5659.5 324 ;
      RECT 5644.5 329 5659.5 344 ;
      RECT 5600 287.5 5615 302.5 ;
      RECT 5580 287.5 5595 302.5 ;
      RECT 5560 287.5 5575 302.5 ;
      RECT 5509.5 361.5 5524.5 376.5 ;
      RECT 5509.5 381.5 5524.5 396.5 ;
      RECT 5509.5 401.5 5524.5 416.5 ;
      RECT 5509.5 451 5524.5 466 ;
      RECT 5509.5 471 5524.5 486 ;
      RECT 5509.5 491 5524.5 506 ;
      RECT 4944.5 119.5 4959.5 134.5 ;
      RECT 4944.5 152 4959.5 167 ;
      RECT 4944.5 697 4959.5 712 ;
      RECT 4944.5 729.5 4959.5 744.5 ;
      RECT 4924.5 119.5 4939.5 134.5 ;
      RECT 4924.5 152 4939.5 167 ;
      RECT 4924.5 697 4939.5 712 ;
      RECT 4924.5 729.5 4939.5 744.5 ;
      RECT 4904.5 119.5 4919.5 134.5 ;
      RECT 4904.5 152 4919.5 167 ;
      RECT 4904.5 697 4919.5 712 ;
      RECT 4904.5 729.5 4919.5 744.5 ;
      RECT 4884.5 119.5 4899.5 134.5 ;
      RECT 4884.5 152 4899.5 167 ;
      RECT 4884.5 697 4899.5 712 ;
      RECT 4884.5 729.5 4899.5 744.5 ;
      RECT 4862.5 343 4877.5 358 ;
      RECT 4862.5 363 4877.5 378 ;
      RECT 4862.5 486 4877.5 501 ;
      RECT 4862.5 506 4877.5 521 ;
      RECT 4842.5 343 4857.5 358 ;
      RECT 4842.5 363 4857.5 378 ;
      RECT 4842.5 486 4857.5 501 ;
      RECT 4842.5 506 4857.5 521 ;
      RECT 4822.5 343 4837.5 358 ;
      RECT 4822.5 363 4837.5 378 ;
      RECT 4822.5 486 4837.5 501 ;
      RECT 4822.5 506 4837.5 521 ;
      RECT 4802.5 343 4817.5 358 ;
      RECT 4802.5 363 4817.5 378 ;
      RECT 4802.5 486 4817.5 501 ;
      RECT 4802.5 506 4817.5 521 ;
      RECT 4750 335.5 4765 350.5 ;
      RECT 4750 513.5 4765 528.5 ;
      RECT 4730 335.5 4745 350.5 ;
      RECT 4730 513.5 4745 528.5 ;
      RECT 4710 335.5 4725 350.5 ;
      RECT 4710 513.5 4725 528.5 ;
      RECT 4705.5 390 4720.5 405 ;
      RECT 4705.5 424.5 4720.5 439.5 ;
      RECT 4705.5 459 4720.5 474 ;
      RECT 4690 335.5 4705 350.5 ;
      RECT 4690 513.5 4705 528.5 ;
      RECT 4685.5 390 4700.5 405 ;
      RECT 4685.5 424.5 4700.5 439.5 ;
      RECT 4685.5 459 4700.5 474 ;
      RECT 4675 182.5 4690 197.5 ;
      RECT 4669.5 666.5 4684.5 681.5 ;
      RECT 4665.5 390 4680.5 405 ;
      RECT 4665.5 424.5 4680.5 439.5 ;
      RECT 4665.5 459 4680.5 474 ;
      RECT 4655 182.5 4670 197.5 ;
      RECT 4649.5 666.5 4664.5 681.5 ;
      RECT 4645.5 390 4660.5 405 ;
      RECT 4645.5 424.5 4660.5 439.5 ;
      RECT 4645.5 459 4660.5 474 ;
      RECT 4635 182.5 4650 197.5 ;
      RECT 4629.5 666.5 4644.5 681.5 ;
      RECT 4615 182.5 4630 197.5 ;
      RECT 4609.5 666.5 4624.5 681.5 ;
      RECT 4493.5 666.5 4508.5 681.5 ;
      RECT 4488.5 182.5 4503.5 197.5 ;
      RECT 4473.5 666.5 4488.5 681.5 ;
      RECT 4468.5 182.5 4483.5 197.5 ;
      RECT 4453.5 666.5 4468.5 681.5 ;
      RECT 4448.5 182.5 4463.5 197.5 ;
      RECT 4433.5 666.5 4448.5 681.5 ;
      RECT 4428.5 182.5 4443.5 197.5 ;
      RECT 4008.5 119.5 4023.5 134.5 ;
      RECT 3988.5 119.5 4003.5 134.5 ;
      RECT 3968.5 119.5 3983.5 134.5 ;
      RECT 3967.5 779 3982.5 794 ;
      RECT 3948.5 119.5 3963.5 134.5 ;
      RECT 3947.5 779 3962.5 794 ;
      RECT 3927.5 779 3942.5 794 ;
      RECT 3907.5 779 3922.5 794 ;
      RECT 3896.5 343 3911.5 358 ;
      RECT 3896.5 363 3911.5 378 ;
      RECT 3896.5 486 3911.5 501 ;
      RECT 3896.5 506 3911.5 521 ;
      RECT 3876.5 343 3891.5 358 ;
      RECT 3876.5 363 3891.5 378 ;
      RECT 3876.5 486 3891.5 501 ;
      RECT 3876.5 506 3891.5 521 ;
      RECT 3868 119.5 3883 134.5 ;
      RECT 3856.5 343 3871.5 358 ;
      RECT 3856.5 363 3871.5 378 ;
      RECT 3856.5 486 3871.5 501 ;
      RECT 3856.5 506 3871.5 521 ;
      RECT 3848 119.5 3863 134.5 ;
      RECT 3836.5 343 3851.5 358 ;
      RECT 3836.5 363 3851.5 378 ;
      RECT 3836.5 486 3851.5 501 ;
      RECT 3836.5 506 3851.5 521 ;
      RECT 3828 119.5 3843 134.5 ;
      RECT 3808 119.5 3823 134.5 ;
      RECT 3784 335.5 3799 350.5 ;
      RECT 3784 513.5 3799 528.5 ;
      RECT 3764 335.5 3779 350.5 ;
      RECT 3764 513.5 3779 528.5 ;
      RECT 3744 335.5 3759 350.5 ;
      RECT 3744 513.5 3759 528.5 ;
      RECT 3739.5 390 3754.5 405 ;
      RECT 3739.5 424.5 3754.5 439.5 ;
      RECT 3739.5 459 3754.5 474 ;
      RECT 3724 335.5 3739 350.5 ;
      RECT 3724 513.5 3739 528.5 ;
      RECT 3719.5 390 3734.5 405 ;
      RECT 3719.5 424.5 3734.5 439.5 ;
      RECT 3719.5 459 3734.5 474 ;
      RECT 3699.5 390 3714.5 405 ;
      RECT 3699.5 424.5 3714.5 439.5 ;
      RECT 3699.5 459 3714.5 474 ;
      RECT 3679.5 390 3694.5 405 ;
      RECT 3679.5 424.5 3694.5 439.5 ;
      RECT 3679.5 459 3694.5 474 ;
      RECT 3658.5 72.5 3673.5 87.5 ;
      RECT 3654.5 155.5 3669.5 170.5 ;
      RECT 3638.5 72.5 3653.5 87.5 ;
      RECT 3634.5 155.5 3649.5 170.5 ;
      RECT 3618.5 72.5 3633.5 87.5 ;
      RECT 3614.5 155.5 3629.5 170.5 ;
      RECT 3609.5 709.5 3624.5 724.5 ;
      RECT 3598.5 72.5 3613.5 87.5 ;
      RECT 3594.5 155.5 3609.5 170.5 ;
      RECT 3589.5 709.5 3604.5 724.5 ;
      RECT 3569.5 709.5 3584.5 724.5 ;
      RECT 3549.5 709.5 3564.5 724.5 ;
      RECT 3547 422 3562 437 ;
      RECT 3547 442 3562 457 ;
      RECT 3547 462 3562 477 ;
      RECT 3530.5 182.5 3545.5 197.5 ;
      RECT 3527 422 3542 437 ;
      RECT 3527 442 3542 457 ;
      RECT 3527 462 3542 477 ;
      RECT 3510.5 182.5 3525.5 197.5 ;
      RECT 3492 287.5 3507 302.5 ;
      RECT 3490.5 182.5 3505.5 197.5 ;
      RECT 3472 287.5 3487 302.5 ;
      RECT 3470.5 182.5 3485.5 197.5 ;
      RECT 3469.5 327.5 3484.5 342.5 ;
      RECT 3469.5 347.5 3484.5 362.5 ;
      RECT 3469.5 367.5 3484.5 382.5 ;
      RECT 3469.5 535.5 3484.5 550.5 ;
      RECT 3469.5 555.5 3484.5 570.5 ;
      RECT 3469.5 575.5 3484.5 590.5 ;
      RECT 3469.5 595.5 3484.5 610.5 ;
      RECT 3452 287.5 3467 302.5 ;
      RECT 3409.5 358.5 3424.5 373.5 ;
      RECT 3409.5 378.5 3424.5 393.5 ;
      RECT 3409.5 398.5 3424.5 413.5 ;
      RECT 3409.5 442.5 3424.5 457.5 ;
      RECT 3409.5 462.5 3424.5 477.5 ;
      RECT 3409.5 482.5 3424.5 497.5 ;
      RECT 3355.5 182.5 3370.5 197.5 ;
      RECT 3335.5 182.5 3350.5 197.5 ;
      RECT 3315.5 182.5 3330.5 197.5 ;
      RECT 3295.5 182.5 3310.5 197.5 ;
      RECT 2844.5 119.5 2859.5 134.5 ;
      RECT 2844.5 152 2859.5 167 ;
      RECT 2826 697 2841 712 ;
      RECT 2826 729.5 2841 744.5 ;
      RECT 2824.5 119.5 2839.5 134.5 ;
      RECT 2824.5 152 2839.5 167 ;
      RECT 2806 697 2821 712 ;
      RECT 2806 729.5 2821 744.5 ;
      RECT 2804.5 119.5 2819.5 134.5 ;
      RECT 2804.5 152 2819.5 167 ;
      RECT 2786 697 2801 712 ;
      RECT 2786 729.5 2801 744.5 ;
      RECT 2784.5 119.5 2799.5 134.5 ;
      RECT 2784.5 152 2799.5 167 ;
      RECT 2766 697 2781 712 ;
      RECT 2766 729.5 2781 744.5 ;
      RECT 2762.5 343 2777.5 358 ;
      RECT 2762.5 363 2777.5 378 ;
      RECT 2762.5 486 2777.5 501 ;
      RECT 2762.5 506 2777.5 521 ;
      RECT 2742.5 343 2757.5 358 ;
      RECT 2742.5 363 2757.5 378 ;
      RECT 2742.5 486 2757.5 501 ;
      RECT 2742.5 506 2757.5 521 ;
      RECT 2722.5 343 2737.5 358 ;
      RECT 2722.5 363 2737.5 378 ;
      RECT 2722.5 486 2737.5 501 ;
      RECT 2722.5 506 2737.5 521 ;
      RECT 2702.5 343 2717.5 358 ;
      RECT 2702.5 363 2717.5 378 ;
      RECT 2702.5 486 2717.5 501 ;
      RECT 2702.5 506 2717.5 521 ;
      RECT 2650 335.5 2665 350.5 ;
      RECT 2650 513.5 2665 528.5 ;
      RECT 2630 335.5 2645 350.5 ;
      RECT 2630 513.5 2645 528.5 ;
      RECT 2610 335.5 2625 350.5 ;
      RECT 2610 513.5 2625 528.5 ;
      RECT 2605.5 390 2620.5 405 ;
      RECT 2605.5 424.5 2620.5 439.5 ;
      RECT 2605.5 459 2620.5 474 ;
      RECT 2590 335.5 2605 350.5 ;
      RECT 2590 513.5 2605 528.5 ;
      RECT 2585.5 390 2600.5 405 ;
      RECT 2585.5 424.5 2600.5 439.5 ;
      RECT 2585.5 459 2600.5 474 ;
      RECT 2579.5 666.5 2594.5 681.5 ;
      RECT 2569.5 182.5 2584.5 197.5 ;
      RECT 2565.5 390 2580.5 405 ;
      RECT 2565.5 424.5 2580.5 439.5 ;
      RECT 2565.5 459 2580.5 474 ;
      RECT 2559.5 666.5 2574.5 681.5 ;
      RECT 2549.5 182.5 2564.5 197.5 ;
      RECT 2545.5 390 2560.5 405 ;
      RECT 2545.5 424.5 2560.5 439.5 ;
      RECT 2545.5 459 2560.5 474 ;
      RECT 2539.5 666.5 2554.5 681.5 ;
      RECT 2529.5 182.5 2544.5 197.5 ;
      RECT 2519.5 666.5 2534.5 681.5 ;
      RECT 2509.5 182.5 2524.5 197.5 ;
      RECT 2393.5 182.5 2408.5 197.5 ;
      RECT 2393.5 666.5 2408.5 681.5 ;
      RECT 2373.5 182.5 2388.5 197.5 ;
      RECT 2373.5 666.5 2388.5 681.5 ;
      RECT 2353.5 182.5 2368.5 197.5 ;
      RECT 2353.5 666.5 2368.5 681.5 ;
      RECT 2333.5 182.5 2348.5 197.5 ;
      RECT 2333.5 666.5 2348.5 681.5 ;
      RECT 1887 130 1902 145 ;
      RECT 1867 130 1882 145 ;
      RECT 1847 130 1862 145 ;
      RECT 1827 130 1842 145 ;
      RECT 1796.5 343 1811.5 358 ;
      RECT 1796.5 363 1811.5 378 ;
      RECT 1796.5 486 1811.5 501 ;
      RECT 1796.5 506 1811.5 521 ;
      RECT 1780 130 1795 145 ;
      RECT 1776.5 343 1791.5 358 ;
      RECT 1776.5 363 1791.5 378 ;
      RECT 1776.5 486 1791.5 501 ;
      RECT 1776.5 506 1791.5 521 ;
      RECT 1760 130 1775 145 ;
      RECT 1756.5 343 1771.5 358 ;
      RECT 1756.5 363 1771.5 378 ;
      RECT 1756.5 486 1771.5 501 ;
      RECT 1756.5 506 1771.5 521 ;
      RECT 1740 130 1755 145 ;
      RECT 1736.5 343 1751.5 358 ;
      RECT 1736.5 363 1751.5 378 ;
      RECT 1736.5 486 1751.5 501 ;
      RECT 1736.5 506 1751.5 521 ;
      RECT 1720 130 1735 145 ;
      RECT 1684 335.5 1699 350.5 ;
      RECT 1684 513.5 1699 528.5 ;
      RECT 1664 335.5 1679 350.5 ;
      RECT 1664 513.5 1679 528.5 ;
      RECT 1644 335.5 1659 350.5 ;
      RECT 1644 513.5 1659 528.5 ;
      RECT 1639.5 390 1654.5 405 ;
      RECT 1639.5 424.5 1654.5 439.5 ;
      RECT 1639.5 459 1654.5 474 ;
      RECT 1624 335.5 1639 350.5 ;
      RECT 1624 513.5 1639 528.5 ;
      RECT 1619.5 390 1634.5 405 ;
      RECT 1619.5 424.5 1634.5 439.5 ;
      RECT 1619.5 459 1634.5 474 ;
      RECT 1599.5 390 1614.5 405 ;
      RECT 1599.5 424.5 1614.5 439.5 ;
      RECT 1599.5 459 1614.5 474 ;
      RECT 1579.5 390 1594.5 405 ;
      RECT 1579.5 424.5 1594.5 439.5 ;
      RECT 1579.5 459 1594.5 474 ;
      RECT 1460 427 1475 442 ;
      RECT 1460 447 1475 462 ;
      RECT 1460 467 1475 482 ;
      RECT 1460 487 1475 502 ;
      RECT 1270 272 1285 287 ;
      RECT 1270 292 1285 307 ;
      RECT 1270 312 1285 327 ;
      RECT 1270 332 1285 347 ;
      RECT 1270 382 1285 397 ;
      RECT 1270 402 1285 417 ;
      RECT 1270 422 1285 437 ;
      RECT 1270 442 1285 457 ;
      RECT 774 99 789 114 ;
      RECT 774 119 789 134 ;
      RECT 770.5 367 785.5 382 ;
      RECT 770.5 387 785.5 402 ;
      RECT 770.5 637 785.5 652 ;
      RECT 770.5 657 785.5 672 ;
      RECT 754 99 769 114 ;
      RECT 754 119 769 134 ;
      RECT 750.5 367 765.5 382 ;
      RECT 750.5 387 765.5 402 ;
      RECT 750.5 637 765.5 652 ;
      RECT 750.5 657 765.5 672 ;
      RECT 734 99 749 114 ;
      RECT 734 119 749 134 ;
      RECT 730.5 367 745.5 382 ;
      RECT 730.5 387 745.5 402 ;
      RECT 730.5 637 745.5 652 ;
      RECT 730.5 657 745.5 672 ;
      RECT 714 99 729 114 ;
      RECT 714 119 729 134 ;
      RECT 710.5 367 725.5 382 ;
      RECT 710.5 387 725.5 402 ;
      RECT 710.5 637 725.5 652 ;
      RECT 710.5 657 725.5 672 ;
      RECT 658 126.5 673 141.5 ;
      RECT 658 394.5 673 409.5 ;
      RECT 658 662.5 673 677.5 ;
      RECT 638 126.5 653 141.5 ;
      RECT 638 394.5 653 409.5 ;
      RECT 638 662.5 653 677.5 ;
      RECT 618 126.5 633 141.5 ;
      RECT 618 394.5 633 409.5 ;
      RECT 618 662.5 633 677.5 ;
      RECT 613.5 37.5 628.5 52.5 ;
      RECT 613.5 72 628.5 87 ;
      RECT 613.5 305.5 628.5 320.5 ;
      RECT 613.5 340 628.5 355 ;
      RECT 613.5 573.5 628.5 588.5 ;
      RECT 613.5 608 628.5 623 ;
      RECT 598 126.5 613 141.5 ;
      RECT 598 394.5 613 409.5 ;
      RECT 598 662.5 613 677.5 ;
      RECT 593.5 37.5 608.5 52.5 ;
      RECT 593.5 72 608.5 87 ;
      RECT 593.5 305.5 608.5 320.5 ;
      RECT 593.5 340 608.5 355 ;
      RECT 593.5 573.5 608.5 588.5 ;
      RECT 593.5 608 608.5 623 ;
      RECT 573.5 37.5 588.5 52.5 ;
      RECT 573.5 72 588.5 87 ;
      RECT 573.5 305.5 588.5 320.5 ;
      RECT 573.5 340 588.5 355 ;
      RECT 573.5 573.5 588.5 588.5 ;
      RECT 573.5 608 588.5 623 ;
      RECT 553.5 37.5 568.5 52.5 ;
      RECT 553.5 72 568.5 87 ;
      RECT 553.5 305.5 568.5 320.5 ;
      RECT 553.5 340 568.5 355 ;
      RECT 553.5 573.5 568.5 588.5 ;
      RECT 553.5 608 568.5 623 ;
      RECT 334.5 829.5 349.5 844.5 ;
      RECT 314.5 829.5 329.5 844.5 ;
      RECT 294.5 829.5 309.5 844.5 ;
      RECT 274.5 829.5 289.5 844.5 ;
      RECT 220.5 709.5 235.5 724.5 ;
      RECT 215.5 441.5 230.5 456.5 ;
      RECT 200.5 709.5 215.5 724.5 ;
      RECT 195.5 441.5 210.5 456.5 ;
      RECT 180.5 709.5 195.5 724.5 ;
      RECT 175.5 441.5 190.5 456.5 ;
      RECT 160.5 709.5 175.5 724.5 ;
      RECT 155.5 441.5 170.5 456.5 ;
      RECT 129.5 709.5 144.5 724.5 ;
      RECT 115.5 441.5 130.5 456.5 ;
      RECT 109.5 709.5 124.5 724.5 ;
      RECT 95.5 441.5 110.5 456.5 ;
      RECT 89.5 709.5 104.5 724.5 ;
      RECT 75.5 441.5 90.5 456.5 ;
      RECT 69.5 709.5 84.5 724.5 ;
      RECT 55.5 441.5 70.5 456.5 ;
    LAYER M2 ;
      RECT 4864 685 4990 752 ;
      RECT 4868.5 112 4976.5 179 ;
      POLYGON 4888 386 4792 386 4792 360 4682 360 4682 325 4888 325 ;
      POLYGON 4888 538 4682 538 4682 504.5 4792 504.5 4792 478 4888 478 ;
      RECT 3794 108 4038.5 146 ;
      POLYGON 4001.5 805.5 3462 805.5 3462 523.5 3492 523.5 3492 767.5 4001.5 767.5 ;
      POLYGON 3922 386 3826 386 3826 359 3716 359 3716 325 3922 325 ;
      POLYGON 3922 538.5 3716 538.5 3716 504 3826 504 3826 478 3922 478 ;
      RECT 3576.5 61.5 3688 177.5 ;
      POLYGON 3518.5 314 3496 314 3496 395 3458 395 3458 314 3440.5 314 3440.5 276.5 3518.5 276.5 ;
      RECT 3398 346.5 3435.5 517 ;
      RECT 2771.5 112 2877.5 179 ;
      RECT 2731.5 685 2866 752 ;
      POLYGON 2788 386 2692 386 2692 360 2582 360 2582 325.5 2788 325.5 ;
      POLYGON 2788 539 2582 539 2582 504.5 2692 504.5 2692 478 2788 478 ;
      RECT 1710.5 118.5 1912 156.5 ;
      POLYGON 1822 386 1726 386 1726 360 1616 360 1616 323.5 1822 323.5 ;
      POLYGON 1822 538.5 1616 538.5 1616 504 1726 504 1726 478 1822 478 ;
      RECT 1258.5 258.5 1296.5 467 ;
      POLYGON 796 149 590 149 590 117 700 117 700 91 796 91 ;
      POLYGON 796 419.5 590 419.5 590 385 700 385 700 359 796 359 ;
      POLYGON 796 687.5 590 687.5 590 653 700 653 700 627 796 627 ;
  END
END DFFD1

MACRO FILL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL1 0 0 ;
  SIZE 10 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 870 10 900 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 10 30 ;
    END
  END VSS
END FILL1

MACRO FILL128
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL128 0 0 ;
  SIZE 1280 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 870 1280 900 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 1280 30 ;
    END
  END VSS
END FILL128

MACRO FILL16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL16 0 0 ;
  SIZE 160 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 870 160 900 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 160 30 ;
    END
  END VSS
END FILL16

MACRO FILL2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL2 0 0 ;
  SIZE 20 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 870 20 900 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 20 30 ;
    END
  END VSS
END FILL2

MACRO FILL32
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL32 0 0 ;
  SIZE 320 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 870 320 900 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 320 30 ;
    END
  END VSS
END FILL32

MACRO FILL4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL4 0 0 ;
  SIZE 40 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 870 40 900 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 40 30 ;
    END
  END VSS
END FILL4

MACRO FILL64
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL64 0 0 ;
  SIZE 640 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 870 640 900 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 640 30 ;
    END
  END VSS
END FILL64

MACRO FILL8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL8 0 0 ;
  SIZE 80 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 870 80 900 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0 80 30 ;
    END
  END VSS
END FILL8

MACRO INVD1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD1 0 0 ;
  SIZE 430 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 430 900 0 900 0 870 90 870 90 580 130 580 130 780 110 780 110 870 318 870 318 780 310 780 310 580 350 580 350 780 342 780 342 870 430 870 ;
    END
  END VDD
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30 590 80 680 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 400 780 360 780 360 580 380 580 380 570 280 570 280 580 300 580 300 780 260 780 260 180 300 180 300 380 280 380 280 410 380 410 380 380 360 380 360 180 400 180 ;
    END
  END OUT
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 178 180 248 270 ;
      LAYER M1 ;
        POLYGON 430 30 350 30 350 380 310 380 310 30 208 30 208 400 170 400 170 300 178 300 178 30 0 30 0 0 430 0 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 190 780 140 780 140 580 160 580 160 570 98 570 98 300 130 300 130 400 122 400 122 410 190 410 ;
    LAYER Via1 ;
      RECT 230 600 240 610 ;
      RECT 230 620 240 630 ;
      RECT 230 640 240 650 ;
      RECT 230 660 240 670 ;
      RECT 228 190 238 200 ;
      RECT 228 210 238 220 ;
      RECT 228 230 238 240 ;
      RECT 228 250 238 260 ;
      RECT 188 190 198 200 ;
      RECT 188 210 198 220 ;
      RECT 188 230 198 240 ;
      RECT 188 250 198 260 ;
      RECT 170 600 180 610 ;
      RECT 170 620 180 630 ;
      RECT 170 640 180 650 ;
      RECT 170 660 180 670 ;
      RECT 48.5 600 58.5 610 ;
      RECT 48.5 620 58.5 630 ;
      RECT 48.5 640 58.5 650 ;
      RECT 48.5 660 58.5 670 ;
    LAYER M2 ;
      RECT 160 590 250 680 ;
  END
END INVD1

MACRO INVD2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD2 0 0 ;
  SIZE 592 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 562 780 522 780 522 580 542 580 542 570 454 570 454 580 462 580 462 780 422 780 422 580 430 580 430 570 342 570 342 580 362 580 362 780 322 780 322 180 362 180 362 380 342 380 342 410 422 410 422 180 462 180 462 380 442 380 442 410 542 410 542 380 522 380 522 180 562 180 ;
    END
  END OUT
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 240 180 310 270 ;
      LAYER M1 ;
        POLYGON 592 30 504 30 504 180 512 180 512 380 472 380 472 180 480 180 480 30 404 30 404 180 412 180 412 380 372 380 372 180 380 180 380 30 270 30 270 400 232 400 232 300 240 300 240 30 104 30 104 300 112 300 112 400 74 400 74 30 0 30 0 0 592 0 ;
    END
  END VSS
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30 590 80 680 ;
    END
  END IN
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 592 900 0 900 0 870 160 870 160 780 152 780 152 580 192 580 192 780 184 780 184 870 380 870 380 780 372 780 372 580 412 580 412 780 404 780 404 870 480 870 480 780 472 780 472 580 512 580 512 780 504 780 504 870 592 870 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      POLYGON 252 780 202 780 202 580 222 580 222 570 122 570 122 580 142 580 142 780 102 780 102 410 160 410 160 400 152 400 152 300 192 300 192 400 184 400 184 410 252 410 ;
    LAYER Via1 ;
      RECT 292 600 302 610 ;
      RECT 292 620 302 630 ;
      RECT 292 640 302 650 ;
      RECT 292 660 302 670 ;
      RECT 290 190 300 200 ;
      RECT 290 210 300 220 ;
      RECT 290 230 300 240 ;
      RECT 290 250 300 260 ;
      RECT 250 190 260 200 ;
      RECT 250 210 260 220 ;
      RECT 250 230 260 240 ;
      RECT 250 250 260 260 ;
      RECT 232 600 242 610 ;
      RECT 232 620 242 630 ;
      RECT 232 640 242 650 ;
      RECT 232 660 242 670 ;
      RECT 48.5 600 58.5 610 ;
      RECT 48.5 620 58.5 630 ;
      RECT 48.5 640 58.5 650 ;
      RECT 48.5 660 58.5 670 ;
    LAYER M2 ;
      RECT 222 590 312 680 ;
  END
END INVD2

MACRO INVD4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD4 0 0 ;
  SIZE 908 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46 590 96 680 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 878 780 838 780 838 580 858 580 858 570 770 570 770 580 778 580 778 780 738 780 738 580 746 580 746 570 670 570 670 580 678 580 678 780 638 780 638 580 646 580 646 570 570 570 570 580 578 580 578 780 538 780 538 580 546 580 546 570 458 570 458 580 478 580 478 780 438 780 438 180 478 180 478 380 458 380 458 410 538 410 538 180 578 180 578 380 558 380 558 410 638 410 638 180 678 180 678 380 658 380 658 410 738 410 738 180 778 180 778 380 758 380 758 410 858 410 858 380 838 380 838 180 878 180 ;
    END
  END OUT
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 356 180 426 270 ;
      LAYER M1 ;
        POLYGON 908 30 820 30 820 180 828 180 828 380 788 380 788 180 796 180 796 30 720 30 720 180 728 180 728 380 688 380 688 180 696 180 696 30 620 30 620 180 628 180 628 380 588 380 588 180 596 180 596 30 520 30 520 180 528 180 528 380 488 380 488 180 496 180 496 30 386 30 386 400 348 400 348 300 356 300 356 30 220 30 220 300 228 300 228 400 188 400 188 300 196 300 196 30 60 30 60 300 68 300 68 400 30 400 30 30 0 30 0 0 908 0 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 908 900 0 900 0 870 176 870 176 780 168 780 168 580 208 580 208 780 200 780 200 870 276 870 276 780 268 780 268 580 308 580 308 780 300 780 300 870 496 870 496 780 488 780 488 580 528 580 528 780 520 780 520 870 596 870 596 780 588 780 588 580 628 580 628 780 620 780 620 870 696 870 696 780 688 780 688 580 728 580 728 780 720 780 720 870 796 870 796 780 788 780 788 580 828 580 828 780 820 780 820 870 908 870 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      POLYGON 368 780 318 780 318 580 338 580 338 570 250 570 250 580 258 580 258 780 218 780 218 580 226 580 226 570 138 570 138 580 158 580 158 780 118 780 118 410 116 410 116 400 108 400 108 300 148 300 148 400 140 400 140 410 276 410 276 400 268 400 268 300 308 300 308 400 300 400 300 410 368 410 ;
    LAYER Via1 ;
      RECT 408 600 418 610 ;
      RECT 408 620 418 630 ;
      RECT 408 640 418 650 ;
      RECT 408 660 418 670 ;
      RECT 406 190 416 200 ;
      RECT 406 210 416 220 ;
      RECT 406 230 416 240 ;
      RECT 406 250 416 260 ;
      RECT 366 190 376 200 ;
      RECT 366 210 376 220 ;
      RECT 366 230 376 240 ;
      RECT 366 250 376 260 ;
      RECT 348 600 358 610 ;
      RECT 348 620 358 630 ;
      RECT 348 640 358 650 ;
      RECT 348 660 358 670 ;
      RECT 64.5 600 74.5 610 ;
      RECT 64.5 620 74.5 630 ;
      RECT 64.5 640 74.5 650 ;
      RECT 64.5 660 74.5 670 ;
    LAYER M2 ;
      RECT 338 590 428 680 ;
  END
END INVD4

MACRO INVD8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD8 0 0 ;
  SIZE 1640 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 1640 900 0 900 0 870 308 870 308 780 300 780 300 580 340 580 340 780 332 780 332 870 408 870 408 780 400 780 400 580 440 580 440 780 432 780 432 870 508 870 508 780 500 780 500 580 540 580 540 780 532 780 532 870 608 870 608 780 600 780 600 580 640 580 640 780 632 780 632 870 828 870 828 780 820 780 820 580 860 580 860 780 852 780 852 870 928 870 928 780 920 780 920 580 960 580 960 780 952 780 952 870 1028 870 1028 780 1020 780 1020 580 1060 580 1060 780 1052 780 1052 870 1128 870 1128 780 1120 780 1120 580 1160 580 1160 780 1152 780 1152 870 1228 870 1228 780 1220 780 1220 580 1260 580 1260 780 1252 780 1252 870 1328 870 1328 780 1320 780 1320 580 1360 580 1360 780 1352 780 1352 870 1428 870 1428 780 1420 780 1420 580 1460 580 1460 780 1452 780 1452 870 1528 870 1528 780 1520 780 1520 580 1560 580 1560 780 1552 780 1552 870 1640 870 ;
    END
  END VDD
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178 590.5 228 680.5 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1610 780 1570 780 1570 580 1590 580 1590 570 1502 570 1502 580 1510 580 1510 780 1470 780 1470 580 1478 580 1478 570 1402 570 1402 580 1410 580 1410 780 1370 780 1370 580 1378 580 1378 570 1302 570 1302 580 1310 580 1310 780 1270 780 1270 580 1278 580 1278 570 1202 570 1202 580 1210 580 1210 780 1170 780 1170 580 1178 580 1178 570 1102 570 1102 580 1110 580 1110 780 1070 780 1070 580 1078 580 1078 570 1002 570 1002 580 1010 580 1010 780 970 780 970 580 978 580 978 570 902 570 902 580 910 580 910 780 870 780 870 580 878 580 878 570 790 570 790 580 810 580 810 780 770 780 770 180 810 180 810 380 790 380 790 410 878 410 878 380 870 380 870 180 910 180 910 380 902 380 902 410 978 410 978 380 970 380 970 180 1010 180 1010 380 1002 380 1002 410 1078 410 1078 380 1070 380 1070 180 1110 180 1110 380 1102 380 1102 410 1178 410 1178 380 1170 380 1170 180 1210 180 1210 380 1202 380 1202 410 1278 410 1278 380 1270 380 1270 180 1310 180 1310 380 1302 380 1302 410 1378 410 1378 380 1370 380 1370 180 1410 180 1410 380 1402 380 1402 410 1478 410 1478 380 1470 380 1470 180 1510 180 1510 380 1502 380 1502 410 1590 410 1590 380 1570 380 1570 180 1610 180 ;
    END
  END OUT
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 688 180 758 270 ;
      LAYER M1 ;
        POLYGON 1640 30 1552 30 1552 180 1560 180 1560 380 1520 380 1520 180 1528 180 1528 30 1452 30 1452 180 1460 180 1460 380 1420 380 1420 180 1428 180 1428 30 1352 30 1352 180 1360 180 1360 380 1320 380 1320 180 1328 180 1328 30 1252 30 1252 180 1260 180 1260 380 1220 380 1220 180 1228 180 1228 30 1152 30 1152 180 1160 180 1160 380 1120 380 1120 180 1128 180 1128 30 1052 30 1052 180 1060 180 1060 380 1020 380 1020 180 1028 180 1028 30 952 30 952 180 960 180 960 380 920 380 920 180 928 180 928 30 852 30 852 180 860 180 860 380 820 380 820 180 828 180 828 30 718 30 718 400 680 400 680 300 688 300 688 30 552 30 552 300 560 300 560 400 520 400 520 300 528 300 528 30 392 30 392 300 400 300 400 400 360 400 360 300 368 300 368 30 232 30 232 300 240 300 240 400 200 400 200 300 208 300 208 30 60 30 60 300 80 300 80 400 30 400 30 30 0 30 0 0 1640 0 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 717.5 570 700 570 700 780 650 780 650 580 670 580 670 570 582 570 582 580 590 580 590 780 550 780 550 580 558 580 558 570 482 570 482 580 490 580 490 780 450 780 450 580 458 580 458 570 382 570 382 580 390 580 390 780 350 780 350 580 358 580 358 570 270 570 270 580 290 580 290 780 250 780 250 570 145.5 570 145.5 410 128 410 128 400 120 400 120 300 160 300 160 400 152 400 152 410 288 410 288 400 280 400 280 300 320 300 320 400 312 400 312 410 448 410 448 400 440 400 440 300 480 300 480 400 472 400 472 410 608 410 608 400 600 400 600 300 640 300 640 400 632 400 632 410 717.5 410 ;
    LAYER Via1 ;
      RECT 740 600 750 610 ;
      RECT 740 620 750 630 ;
      RECT 740 640 750 650 ;
      RECT 740 660 750 670 ;
      RECT 738 190 748 200 ;
      RECT 738 210 748 220 ;
      RECT 738 230 748 240 ;
      RECT 738 250 748 260 ;
      RECT 698 190 708 200 ;
      RECT 698 210 708 220 ;
      RECT 698 230 708 240 ;
      RECT 698 250 708 260 ;
      RECT 680 600 690 610 ;
      RECT 680 620 690 630 ;
      RECT 680 640 690 650 ;
      RECT 680 660 690 670 ;
      RECT 196.5 600.5 206.5 610.5 ;
      RECT 196.5 620.5 206.5 630.5 ;
      RECT 196.5 640.5 206.5 650.5 ;
      RECT 196.5 660.5 206.5 670.5 ;
    LAYER M2 ;
      RECT 670 590 760 680 ;
  END
END INVD8

MACRO NAND2D1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2D1 0 0 ;
  SIZE 610 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 520 830 490 830 490 581.7 440 581.7 440 830 410 830 410 538.9 200 538.9 200 830 170 830 170 581.7 120 581.7 120 830 90 830 90 522.8 371.4 522.8 371.4 256.6 401.4 256.6 401.4 522.8 451.4 522.8 451.4 256.6 481.4 256.6 481.4 522.8 520 522.8 ;
    END
  END OUT
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 276.1 418.4 204.1 418.4 204.1 329.3 132.1 329.3 132.1 283.3 276.1 283.3 ;
      LAYER M1 ;
        POLYGON 610 30 521.4 30 521.4 456.6 491.4 456.6 491.4 239.3 441.4 239.3 441.4 456.6 411.4 456.6 411.4 239.3 361.4 239.3 361.4 456.6 179.7 456.6 179.7 472.4 150 472.4 150 372.4 331.4 372.4 331.4 30 0 30 0 0 610 0 ;
    END
  END VSS
  PIN IN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 565 612 595 702 ;
    END
  END IN2
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 610 900 0 900 0 870 60 870 60 630 80 630 80 870 130 870 130 630 160 630 160 870 210 870 210 630 240 630 240 870 290 870 290 630 320 630 320 870 370 870 370 630 400 630 400 870 450 870 450 630 480 630 480 870 530 870 530 630 550 630 550 870 610 870 ;
    END
  END VDD
  PIN IN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15 612 45 702 ;
    END
  END IN1
  OBS
    LAYER M1 ;
      POLYGON 360 830 330 830 330 583.1 280 583.1 280 830 250 830 250 558.7 360 558.7 ;
      POLYGON 180.5 503.9 121.5 503.9 121.5 486.9 120 486.9 120 372.4 140 372.4 140 483.9 180.5 483.9 ;
    LAYER Via1 ;
      RECT 575 622 585 632 ;
      RECT 575 642 585 652 ;
      RECT 575 662 585 672 ;
      RECT 575 682 585 692 ;
      RECT 318.9 568.1 326.9 576.1 ;
      RECT 317.1 489.9 325.1 497.9 ;
      RECT 305.9 568.1 313.9 576.1 ;
      RECT 304.1 489.9 312.1 497.9 ;
      RECT 292.9 568.1 300.9 576.1 ;
      RECT 291.1 489.9 299.1 497.9 ;
      RECT 279.9 568.1 287.9 576.1 ;
      RECT 278.1 489.9 286.1 497.9 ;
      RECT 262.1 378.4 270.1 386.4 ;
      RECT 262.1 391.4 270.1 399.4 ;
      RECT 262.1 404.4 270.1 412.4 ;
      RECT 249.1 378.4 257.1 386.4 ;
      RECT 249.1 391.4 257.1 399.4 ;
      RECT 249.1 404.4 257.1 412.4 ;
      RECT 236.1 378.4 244.1 386.4 ;
      RECT 236.1 391.4 244.1 399.4 ;
      RECT 236.1 404.4 244.1 412.4 ;
      RECT 223.1 378.4 231.1 386.4 ;
      RECT 223.1 391.4 231.1 399.4 ;
      RECT 223.1 404.4 231.1 412.4 ;
      RECT 210.1 378.4 218.1 386.4 ;
      RECT 210.1 391.4 218.1 399.4 ;
      RECT 210.1 404.4 218.1 412.4 ;
      RECT 190.1 289.3 198.1 297.3 ;
      RECT 190.1 302.3 198.1 310.3 ;
      RECT 190.1 315.3 198.1 323.3 ;
      RECT 177.1 289.3 185.1 297.3 ;
      RECT 177.1 302.3 185.1 310.3 ;
      RECT 177.1 315.3 185.1 323.3 ;
      RECT 166.5 489.9 174.5 497.9 ;
      RECT 164.1 289.3 172.1 297.3 ;
      RECT 164.1 302.3 172.1 310.3 ;
      RECT 164.1 315.3 172.1 323.3 ;
      RECT 153.5 489.9 161.5 497.9 ;
      RECT 151.1 289.3 159.1 297.3 ;
      RECT 151.1 302.3 159.1 310.3 ;
      RECT 151.1 315.3 159.1 323.3 ;
      RECT 140.5 489.9 148.5 497.9 ;
      RECT 138.1 289.3 146.1 297.3 ;
      RECT 138.1 302.3 146.1 310.3 ;
      RECT 138.1 315.3 146.1 323.3 ;
      RECT 127.5 489.9 135.5 497.9 ;
      RECT 25 622 35 632 ;
      RECT 25 642 35 652 ;
      RECT 25 662 35 672 ;
      RECT 25 682 35 692 ;
    LAYER M2 ;
      POLYGON 344.4 584.2 261.1 584.2 261.1 505.2 117 505.2 117 483.4 344.4 483.4 ;
  END
END NAND2D1

MACRO NAND2D2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2D2 0 0 ;
  SIZE 610 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN IN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 565 612 595 702 ;
    END
  END IN2
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 183.5 236 163.5 236 163.5 141.2 101.2 141.2 101.2 121.2 183.5 121.2 ;
      LAYER M1 ;
        POLYGON 610 30 574.6 30 574.6 243.6 544.6 243.6 544.6 30 494.6 30 494.6 243.6 464.6 243.6 464.6 30 414.6 30 414.6 243.6 384.6 243.6 384.6 30 334.6 30 334.6 243.6 304.6 243.6 304.6 30 254.6 30 254.6 243.6 170 243.6 170 272.4 150 272.4 150 160 100 160 100 272.4 80 272.4 80 145 170 145 170 172.4 224.6 172.4 224.6 30 0 30 0 0 610 0 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 610 900 0 900 0 870 60 870 60 430 80 430 80 870 130 870 130 430 160 430 160 870 210 870 210 430 240 430 240 870 290 870 290 430 320 430 320 870 370 870 370 430 400 430 400 870 450 870 450 430 480 430 480 870 530 870 530 430 550 430 550 870 610 870 ;
    END
  END VDD
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 534.6 356 520 356 520 830 490 830 490 381.7 440 381.7 440 830 410 830 410 338.9 200 338.9 200 830 170 830 170 381.7 120 381.7 120 830 90 830 90 322.8 504.6 322.8 504.6 273.3 264.6 273.3 264.6 43.6 294.6 43.6 294.6 243.6 294.7 243.6 294.7 258.6 344.6 258.6 344.6 43.6 374.6 43.6 374.6 258.6 424.6 258.6 424.6 43.6 454.6 43.6 454.6 243.6 454.7 243.6 454.7 258.6 504.6 258.6 504.6 43.6 534.6 43.6 ;
    END
  END OUT
  PIN IN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15 612 45 702 ;
    END
  END IN1
  OBS
    LAYER M1 ;
      POLYGON 360 830 330 830 330 383.1 280 383.1 280 830 250 830 250 358.7 360 358.7 ;
      POLYGON 180.5 303.9 80 303.9 80 283.9 110 283.9 110 172.4 140 172.4 140 283.9 180.5 283.9 ;
    LAYER Via1 ;
      RECT 575 622 585 632 ;
      RECT 575 642 585 652 ;
      RECT 575 662 585 672 ;
      RECT 575 682 585 692 ;
      RECT 318.9 368.1 326.9 376.1 ;
      RECT 317.1 289.9 325.1 297.9 ;
      RECT 305.9 368.1 313.9 376.1 ;
      RECT 304.1 289.9 312.1 297.9 ;
      RECT 292.9 368.1 300.9 376.1 ;
      RECT 291.1 289.9 299.1 297.9 ;
      RECT 279.9 368.1 287.9 376.1 ;
      RECT 278.1 289.9 286.1 297.9 ;
      RECT 169.5 183 177.5 191 ;
      RECT 169.5 196 177.5 204 ;
      RECT 169.5 209 177.5 217 ;
      RECT 169.5 222 177.5 230 ;
      RECT 166.5 289.9 174.5 297.9 ;
      RECT 153.5 289.9 161.5 297.9 ;
      RECT 146.2 127.2 154.2 135.2 ;
      RECT 140.5 289.9 148.5 297.9 ;
      RECT 133.2 127.2 141.2 135.2 ;
      RECT 127.5 289.9 135.5 297.9 ;
      RECT 120.2 127.2 128.2 135.2 ;
      RECT 107.2 127.2 115.2 135.2 ;
      RECT 25 622 35 632 ;
      RECT 25 642 35 652 ;
      RECT 25 662 35 672 ;
      RECT 25 682 35 692 ;
    LAYER M2 ;
      POLYGON 344.4 384.2 261.1 384.2 261.1 305.2 117 305.2 117 283.4 344.4 283.4 ;
  END
END NAND2D2

MACRO NAND2D4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2D4 0 0 ;
  SIZE 1090 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN IN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1045 612 1075 702 ;
    END
  END IN2
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 1090 900 0 900 0 870 60 870 60 430 80 430 80 870 130 870 130 430 160 430 160 870 210 870 210 430 240 430 240 870 290 870 290 430 320 430 320 870 370 870 370 430 400 430 400 870 450 870 450 430 480 430 480 870 530 870 530 430 560 430 560 870 610 870 610 430 640 430 640 870 690 870 690 430 720 430 720 870 770 870 770 430 800 430 800 870 850 870 850 430 880 430 880 870 930 870 930 430 960 430 960 870 1010 870 1010 430 1030 430 1030 870 1090 870 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 328.9 236 308.9 236 308.9 141.2 244.5 141.2 244.5 121.2 328.9 121.2 ;
      LAYER M1 ;
        POLYGON 1090 30 1030 30 1030 243.6 1010 243.6 1010 30 960 30 960 243.6 930 243.6 930 30 880 30 880 243.6 850 243.6 850 30 800 30 800 243.6 770 243.6 770 30 720 30 720 243.6 690 243.6 690 30 640 30 640 243.6 610 243.6 610 30 560 30 560 243.6 530 243.6 530 30 480 30 480 243.6 450 243.6 450 30 400 30 400 243.6 310 243.6 310 272.4 295.4 272.4 295.4 159.9 245.4 159.9 245.4 272.4 215.4 272.4 215.4 159.9 165.4 159.9 165.4 272.4 145.4 272.4 145.4 145 310 145 310 172.4 370 172.4 370 30 0 30 0 0 1090 0 ;
    END
  END VSS
  PIN IN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15 613 45 703 ;
    END
  END IN1
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1000 273.3 680 273.3 680 322.8 1000 322.8 1000 830 970 830 970 338.9 920 338.9 920 830 890 830 890 338.9 840 338.9 840 830 810 830 810 338.9 760 338.9 760 830 730 830 730 338.9 360 338.9 360 830 330 830 330 338.9 280 338.9 280 830 250 830 250 338.9 200 338.9 200 830 170 830 170 338.9 120 338.9 120 830 90 830 90 322.8 650 322.8 650 273.3 410 273.3 410 43.6 440 43.6 440 243.6 440.1 243.6 440.1 258.6 490 258.6 490 43.6 520 43.6 520 258.6 570 258.6 570 43.6 600 43.6 600 243.6 600.1 243.6 600.1 258.6 650 258.6 650 43.6 680 43.6 680 258.6 730 258.6 730 43.6 760 43.6 760 243.6 760.1 243.6 760.1 258.6 810 258.6 810 43.6 840 43.6 840 258.6 890 258.6 890 43.6 920 43.6 920 243.6 920.1 243.6 920.1 258.6 970 258.6 970 43.6 1000 43.6 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      POLYGON 680 830 650 830 650 383.1 600 383.1 600 830 570 830 570 383.1 520 383.1 520 830 490 830 490 383.1 440 383.1 440 830 410 830 410 358.7 680 358.7 ;
      POLYGON 325.9 303.9 155.4 303.9 155.4 283.9 175.4 283.9 175.4 172.4 205.4 172.4 205.4 272.4 205.5 272.4 205.5 283.9 255.4 283.9 255.4 172.4 285.4 172.4 285.4 283.9 325.9 283.9 ;
    LAYER Via1 ;
      RECT 1055 622 1065 632 ;
      RECT 1055 642 1065 652 ;
      RECT 1055 662 1065 672 ;
      RECT 1055 682 1065 692 ;
      RECT 464.3 368.1 472.3 376.1 ;
      RECT 462.5 289.9 470.5 297.9 ;
      RECT 451.3 368.1 459.3 376.1 ;
      RECT 449.5 289.9 457.5 297.9 ;
      RECT 438.3 368.1 446.3 376.1 ;
      RECT 436.5 289.9 444.5 297.9 ;
      RECT 425.3 368.1 433.3 376.1 ;
      RECT 423.5 289.9 431.5 297.9 ;
      RECT 314.9 183 322.9 191 ;
      RECT 314.9 196 322.9 204 ;
      RECT 314.9 209 322.9 217 ;
      RECT 314.9 222 322.9 230 ;
      RECT 311.9 289.9 319.9 297.9 ;
      RECT 298.9 289.9 306.9 297.9 ;
      RECT 289.5 127.2 297.5 135.2 ;
      RECT 285.9 289.9 293.9 297.9 ;
      RECT 276.5 127.2 284.5 135.2 ;
      RECT 272.9 289.9 280.9 297.9 ;
      RECT 263.5 127.2 271.5 135.2 ;
      RECT 250.5 127.2 258.5 135.2 ;
      RECT 25 623 35 633 ;
      RECT 25 643 35 653 ;
      RECT 25 663 35 673 ;
      RECT 25 683 35 693 ;
    LAYER M2 ;
      POLYGON 489.8 384.2 406.5 384.2 406.5 305.2 262.4 305.2 262.4 283.4 489.8 283.4 ;
  END
END NAND2D4

MACRO NAND2D8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2D8 0 0 ;
  SIZE 2050 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 2050 900 0 900 0 870 60 870 60 430 80 430 80 870 130 870 130 430 160 430 160 870 210 870 210 430 240 430 240 870 290 870 290 430 320 430 320 870 370 870 370 430 400 430 400 870 450 870 450 430 480 430 480 870 530 870 530 430 560 430 560 870 610 870 610 430 640 430 640 870 690 870 690 430 720 430 720 870 770 870 770 430 800 430 800 870 850 870 850 430 880 430 880 870 930 870 930 430 960 430 960 870 1010 870 1010 430 1040 430 1040 870 1090 870 1090 430 1120 430 1120 870 1170 870 1170 430 1200 430 1200 870 1250 870 1250 430 1280 430 1280 870 1330 870 1330 430 1360 430 1360 870 1410 870 1410 430 1440 430 1440 870 1490 870 1490 430 1520 430 1520 870 1570 870 1570 430 1600 430 1600 870 1650 870 1650 430 1680 430 1680 870 1730 870 1730 430 1760 430 1760 870 1810 870 1810 430 1840 430 1840 870 1890 870 1890 430 1920 430 1920 870 1970 870 1970 430 1990 430 1990 870 2050 870 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 648.9 236 628.9 236 628.9 141.2 564.5 141.2 564.5 121.2 648.9 121.2 ;
      LAYER M1 ;
        POLYGON 2050 30 1990 30 1990 243.6 1970 243.6 1970 30 1920 30 1920 243.6 1890 243.6 1890 30 1840 30 1840 243.6 1810 243.6 1810 30 1760 30 1760 243.6 1730 243.6 1730 30 1680 30 1680 243.6 1650 243.6 1650 30 1600 30 1600 243.6 1570 243.6 1570 30 1520 30 1520 243.6 1490 243.6 1490 30 1440 30 1440 243.6 1410 243.6 1410 30 1360 30 1360 243.6 1330 243.6 1330 30 1280 30 1280 243.6 1250 243.6 1250 30 1200 30 1200 243.6 1170 243.6 1170 30 1120 30 1120 243.6 1090 243.6 1090 30 1040 30 1040 243.6 1010 243.6 1010 30 960 30 960 243.6 930 243.6 930 30 880 30 880 243.6 850 243.6 850 30 800 30 800 243.6 770 243.6 770 30 720 30 720 243.6 635.4 243.6 635.4 272.4 615.4 272.4 615.4 159.9 565.4 159.9 565.4 272.4 535.4 272.4 535.4 159.9 485.4 159.9 485.4 272.4 455.4 272.4 455.4 159.9 405.4 159.9 405.4 272.4 375.4 272.4 375.4 159.9 325.4 159.9 325.4 272.4 309.4 272.4 309.4 144.5 635.4 144.5 635.4 172.4 690 172.4 690 30 0 30 0 0 2050 0 ;
    END
  END VSS
  PIN IN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2005 612 2035 702 ;
    END
  END IN2
  PIN IN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.5 612 44.5 702 ;
    END
  END IN1
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1960 273.3 1000 273.3 1000 322.8 1960 322.8 1960 830 1930 830 1930 338.9 1880 338.9 1880 830 1850 830 1850 338.9 1800 338.9 1800 830 1770 830 1770 338.9 1720 338.9 1720 830 1690 830 1690 338.9 1640 338.9 1640 830 1610 830 1610 338.9 1560 338.9 1560 830 1530 830 1530 338.9 1480 338.9 1480 830 1450 830 1450 338.9 1400 338.9 1400 830 1370 830 1370 338.9 680 338.9 680 830 650 830 650 338.9 600 338.9 600 830 570 830 570 338.9 520 338.9 520 830 490 830 490 338.9 440 338.9 440 830 410 830 410 338.9 360 338.9 360 830 330 830 330 338.9 280 338.9 280 830 250 830 250 338.9 200 338.9 200 830 170 830 170 338.9 120 338.9 120 830 90 830 90 322.8 970 322.8 970 273.3 730 273.3 730 43.6 760 43.6 760 243.6 760.1 243.6 760.1 258.6 810 258.6 810 43.6 840 43.6 840 258.6 890 258.6 890 43.6 920 43.6 920 243.6 920.1 243.6 920.1 258.6 970 258.6 970 43.6 1000 43.6 1000 258.6 1050 258.6 1050 43.6 1080 43.6 1080 243.6 1080.1 243.6 1080.1 258.6 1130 258.6 1130 43.6 1160 43.6 1160 258.6 1210 258.6 1210 43.6 1240 43.6 1240 243.6 1240.1 243.6 1240.1 258.6 1290 258.6 1290 43.6 1320 43.6 1320 258.6 1370 258.6 1370 43.6 1400 43.6 1400 243.6 1400.1 243.6 1400.1 258.6 1450 258.6 1450 43.6 1480 43.6 1480 258.6 1530 258.6 1530 43.6 1560 43.6 1560 243.6 1560.1 243.6 1560.1 258.6 1610 258.6 1610 43.6 1640 43.6 1640 258.6 1690 258.6 1690 43.6 1720 43.6 1720 243.6 1720.1 243.6 1720.1 258.6 1770 258.6 1770 43.6 1800 43.6 1800 258.6 1850 258.6 1850 43.6 1880 43.6 1880 243.6 1880.1 243.6 1880.1 258.6 1930 258.6 1930 43.6 1960 43.6 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      POLYGON 1320 830 1290 830 1290 383.1 1240 383.1 1240 830 1210 830 1210 383.1 1160 383.1 1160 830 1130 830 1130 383.1 1080 383.1 1080 830 1050 830 1050 383.1 1000 383.1 1000 830 970 830 970 383.1 920 383.1 920 830 890 830 890 383.1 840 383.1 840 830 810 830 810 383.1 760 383.1 760 830 730 830 730 358.7 1320 358.7 ;
      POLYGON 645.9 303.9 309.4 303.9 309.4 283.9 335.4 283.9 335.4 172.4 365.4 172.4 365.4 283.9 415.4 283.9 415.4 172.4 445.4 172.4 445.4 283.9 495.4 283.9 495.4 172.4 525.4 172.4 525.4 283.9 575.4 283.9 575.4 172.4 605.4 172.4 605.4 283.9 645.9 283.9 ;
    LAYER Via1 ;
      RECT 2015 622 2025 632 ;
      RECT 2015 642 2025 652 ;
      RECT 2015 662 2025 672 ;
      RECT 2015 682 2025 692 ;
      RECT 784.3 368.1 792.3 376.1 ;
      RECT 782.5 289.9 790.5 297.9 ;
      RECT 771.3 368.1 779.3 376.1 ;
      RECT 769.5 289.9 777.5 297.9 ;
      RECT 758.3 368.1 766.3 376.1 ;
      RECT 756.5 289.9 764.5 297.9 ;
      RECT 745.3 368.1 753.3 376.1 ;
      RECT 743.5 289.9 751.5 297.9 ;
      RECT 634.9 183 642.9 191 ;
      RECT 634.9 196 642.9 204 ;
      RECT 634.9 209 642.9 217 ;
      RECT 634.9 222 642.9 230 ;
      RECT 631.9 289.9 639.9 297.9 ;
      RECT 618.9 289.9 626.9 297.9 ;
      RECT 609.5 127.2 617.5 135.2 ;
      RECT 605.9 289.9 613.9 297.9 ;
      RECT 596.5 127.2 604.5 135.2 ;
      RECT 592.9 289.9 600.9 297.9 ;
      RECT 583.5 127.2 591.5 135.2 ;
      RECT 570.5 127.2 578.5 135.2 ;
      RECT 24.5 622 34.5 632 ;
      RECT 24.5 642 34.5 652 ;
      RECT 24.5 662 34.5 672 ;
      RECT 24.5 682 34.5 692 ;
    LAYER M2 ;
      POLYGON 809.8 384.2 726.5 384.2 726.5 305.2 582.4 305.2 582.4 283.4 809.8 283.4 ;
  END
END NAND2D8

MACRO NOR2D1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2D1 0 0 ;
  SIZE 520 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 520 900 0 900 0 870 110 870 110 630 140 630 140 870 190 870 190 630 220 630 220 870 340 870 340 630 370 630 370 870 420 870 420 630 450 630 450 870 520 870 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 200 70 270 150 ;
      LAYER M1 ;
        POLYGON 520 30 490 30 490 100 455 100 455 120 355 120 355 100 190 100 190 160 90 160 90 30 0 30 0 0 520 0 ;
    END
  END VSS
  PIN IN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20 292 50 382 ;
    END
  END IN2
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 490 270 450 270 450 510 420 510 420 270 370 270 370 510 340 510 340 270 320 270 320 150 355 150 355 130 455 130 455 150 490 150 ;
    END
  END OUT
  PIN IN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20 612 50 702 ;
    END
  END IN1
  OBS
    LAYER M1 ;
      POLYGON 490 830 460 830 460 590 410 590 410 830 380 830 380 590 330 590 330 830 300 830 300 310 330 310 330 550 380 550 380 310 410 310 410 550 460 550 460 310 490 310 ;
      POLYGON 260 830 230 830 230 590 180 590 180 830 150 830 150 590 100 590 100 830 70 830 70 310 100 310 100 550 150 550 150 310 180 310 180 550 230 550 230 310 260 310 ;
      POLYGON 220 510 190 510 190 270 140 270 140 510 110 510 110 270 90 270 90 170 190 170 190 190 220 190 ;
    LAYER Via1 ;
      RECT 290 240 300 250 ;
      RECT 270 240 280 250 ;
      RECT 250 80 260 90 ;
      RECT 250 130 260 140 ;
      RECT 250 240 260 250 ;
      RECT 230 80 240 90 ;
      RECT 230 130 240 140 ;
      RECT 210 80 220 90 ;
      RECT 210 130 220 140 ;
      RECT 200 240 210 250 ;
      RECT 180 240 190 250 ;
      RECT 160 240 170 250 ;
      RECT 30 302 40 312 ;
      RECT 30 322 40 332 ;
      RECT 30 342 40 352 ;
      RECT 30 362 40 372 ;
      RECT 30 622 40 632 ;
      RECT 30 642 40 652 ;
      RECT 30 662 40 672 ;
      RECT 30 682 40 692 ;
    LAYER M2 ;
      RECT 150 230 310 260 ;
  END
END NOR2D1

MACRO NOR2D2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2D2 0 0 ;
  SIZE 840 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 810 270 770 270 770 510 740 510 740 270 690 270 690 510 660 510 660 270 610 270 610 510 580 510 580 270 530 270 530 510 500 510 500 150 555 150 555 130 755 130 755 150 810 150 ;
    END
  END OUT
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 840 900 0 900 0 870 110 870 110 630 140 630 140 870 190 870 190 630 220 630 220 870 270 870 270 630 300 630 300 870 350 870 350 630 380 630 380 870 500 870 500 630 530 630 530 870 580 870 580 630 610 630 610 870 660 870 660 630 690 630 690 870 740 870 740 630 770 630 770 870 840 870 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 300 70 370 150 ;
      LAYER M1 ;
        POLYGON 840 30 810 30 810 100 755 100 755 120 555 120 555 100 290 100 290 160 90 160 90 30 0 30 0 0 840 0 ;
    END
  END VSS
  PIN IN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20 292 50 382 ;
    END
  END IN2
  PIN IN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.5 612 50.5 702 ;
    END
  END IN1
  OBS
    LAYER M1 ;
      POLYGON 810 830 780 830 780 590 730 590 730 830 700 830 700 590 650 590 650 830 620 830 620 590 570 590 570 830 540 830 540 590 490 590 490 830 460 830 460 310 490 310 490 550 540 550 540 310 570 310 570 550 620 550 620 310 650 310 650 550 700 550 700 310 730 310 730 550 780 550 780 310 810 310 ;
      POLYGON 420 830 390 830 390 590 340 590 340 830 310 830 310 590 260 590 260 830 230 830 230 590 180 590 180 830 150 830 150 590 100 590 100 830 70 830 70 310 100 310 100 550 150 550 150 310 180 310 180 550 230 550 230 310 260 310 260 550 310 550 310 310 340 310 340 550 390 550 390 310 420 310 ;
      POLYGON 380 510 350 510 350 270 300 270 300 510 270 510 270 270 220 270 220 510 190 510 190 270 140 270 140 510 110 510 110 270 90 270 90 170 290 170 290 190 380 190 ;
    LAYER Via1 ;
      RECT 450 240 460 250 ;
      RECT 430 240 440 250 ;
      RECT 410 240 420 250 ;
      RECT 360 240 370 250 ;
      RECT 350 80 360 90 ;
      RECT 350 130 360 140 ;
      RECT 340 240 350 250 ;
      RECT 330 80 340 90 ;
      RECT 330 130 340 140 ;
      RECT 320 240 330 250 ;
      RECT 310 80 320 90 ;
      RECT 310 130 320 140 ;
      RECT 30.5 622 40.5 632 ;
      RECT 30.5 642 40.5 652 ;
      RECT 30.5 662 40.5 672 ;
      RECT 30.5 682 40.5 692 ;
      RECT 30 302 40 312 ;
      RECT 30 322 40 332 ;
      RECT 30 342 40 352 ;
      RECT 30 362 40 372 ;
    LAYER M2 ;
      RECT 310 230 470 260 ;
  END
END NOR2D2

MACRO NOR2D4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2D4 0 0 ;
  SIZE 1480 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 1480 900 0 900 0 870 110 870 110 630 140 630 140 870 190 870 190 630 220 630 220 870 270 870 270 630 300 630 300 870 350 870 350 630 380 630 380 870 430 870 430 630 460 630 460 870 510 870 510 630 540 630 540 870 590 870 590 630 620 630 620 870 670 870 670 630 700 630 700 870 820 870 820 630 850 630 850 870 900 870 900 630 930 630 930 870 980 870 980 630 1010 630 1010 870 1060 870 1060 630 1090 630 1090 870 1140 870 1140 630 1170 630 1170 870 1220 870 1220 630 1250 630 1250 870 1300 870 1300 630 1330 630 1330 870 1380 870 1380 630 1410 630 1410 870 1480 870 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 500 70 570 150 ;
      LAYER M1 ;
        POLYGON 1480 30 1450 30 1450 100 1335 100 1335 120 935 120 935 100 490 100 490 160 90 160 90 30 0 30 0 0 1480 0 ;
    END
  END VSS
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1450 270 1410 270 1410 510 1380 510 1380 270 1330 270 1330 510 1300 510 1300 270 1250 270 1250 510 1220 510 1220 270 1170 270 1170 510 1140 510 1140 270 1090 270 1090 510 1060 510 1060 270 1010 270 1010 510 980 510 980 270 930 270 930 510 900 510 900 270 850 270 850 510 820 510 820 150 935 150 935 130 1335 130 1335 150 1450 150 ;
    END
  END OUT
  PIN IN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20 292 50 382 ;
    END
  END IN2
  PIN IN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20 612 50 702 ;
    END
  END IN1
  OBS
    LAYER M1 ;
      POLYGON 1450 830 1420 830 1420 590 1370 590 1370 830 1340 830 1340 590 1290 590 1290 830 1260 830 1260 590 1210 590 1210 830 1180 830 1180 590 1130 590 1130 830 1100 830 1100 590 1050 590 1050 830 1020 830 1020 590 970 590 970 830 940 830 940 590 890 590 890 830 860 830 860 590 810 590 810 830 780 830 780 310 810 310 810 550 860 550 860 310 890 310 890 550 940 550 940 310 970 310 970 550 1020 550 1020 310 1050 310 1050 550 1100 550 1100 310 1130 310 1130 550 1180 550 1180 310 1210 310 1210 550 1260 550 1260 310 1290 310 1290 550 1340 550 1340 310 1370 310 1370 550 1420 550 1420 310 1450 310 ;
      POLYGON 740 830 710 830 710 590 660 590 660 830 630 830 630 590 580 590 580 830 550 830 550 590 500 590 500 830 470 830 470 590 420 590 420 830 390 830 390 590 340 590 340 830 310 830 310 590 260 590 260 830 230 830 230 590 180 590 180 830 150 830 150 590 100 590 100 830 70 830 70 310 100 310 100 550 150 550 150 310 180 310 180 550 230 550 230 310 260 310 260 550 310 550 310 310 340 310 340 550 390 550 390 310 420 310 420 550 470 550 470 310 500 310 500 550 550 550 550 310 580 310 580 550 630 550 630 310 660 310 660 550 710 550 710 310 740 310 ;
      POLYGON 700 510 670 510 670 270 620 270 620 510 590 510 590 270 540 270 540 510 510 510 510 270 460 270 460 510 430 510 430 270 380 270 380 510 350 510 350 270 300 270 300 510 270 510 270 270 220 270 220 510 190 510 190 270 140 270 140 510 110 510 110 270 90 270 90 170 490 170 490 190 700 190 ;
    LAYER Via1 ;
      RECT 770 240 780 250 ;
      RECT 750 240 760 250 ;
      RECT 730 240 740 250 ;
      RECT 680 240 690 250 ;
      RECT 660 240 670 250 ;
      RECT 640 240 650 250 ;
      RECT 550 80 560 90 ;
      RECT 550 130 560 140 ;
      RECT 530 80 540 90 ;
      RECT 530 130 540 140 ;
      RECT 510 80 520 90 ;
      RECT 510 130 520 140 ;
      RECT 30 302 40 312 ;
      RECT 30 322 40 332 ;
      RECT 30 342 40 352 ;
      RECT 30 362 40 372 ;
      RECT 30 622 40 632 ;
      RECT 30 642 40 652 ;
      RECT 30 662 40 672 ;
      RECT 30 682 40 692 ;
    LAYER M2 ;
      RECT 630 230 790 260 ;
  END
END NOR2D4

MACRO NOR2D8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2D8 0 0 ;
  SIZE 2760 BY 900 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 2760 900 0 900 0 870 110 870 110 630 140 630 140 870 190 870 190 630 220 630 220 870 270 870 270 630 300 630 300 870 350 870 350 630 380 630 380 870 430 870 430 630 460 630 460 870 510 870 510 630 540 630 540 870 590 870 590 630 620 630 620 870 670 870 670 630 700 630 700 870 750 870 750 630 780 630 780 870 830 870 830 630 860 630 860 870 910 870 910 630 940 630 940 870 990 870 990 630 1020 630 1020 870 1070 870 1070 630 1100 630 1100 870 1150 870 1150 630 1180 630 1180 870 1230 870 1230 630 1260 630 1260 870 1310 870 1310 630 1340 630 1340 870 1460 870 1460 630 1490 630 1490 870 1540 870 1540 630 1570 630 1570 870 1620 870 1620 630 1650 630 1650 870 1700 870 1700 630 1730 630 1730 870 1780 870 1780 630 1810 630 1810 870 1860 870 1860 630 1890 630 1890 870 1940 870 1940 630 1970 630 1970 870 2020 870 2020 630 2050 630 2050 870 2100 870 2100 630 2130 630 2130 870 2180 870 2180 630 2210 630 2210 870 2260 870 2260 630 2290 630 2290 870 2340 870 2340 630 2370 630 2370 870 2420 870 2420 630 2450 630 2450 870 2500 870 2500 630 2530 630 2530 870 2580 870 2580 630 2610 630 2610 870 2660 870 2660 630 2690 630 2690 870 2760 870 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 900 70 970 150 ;
      LAYER M1 ;
        POLYGON 2760 30 2730 30 2730 100 2495 100 2495 120 1695 120 1695 100 890 100 890 160 90 160 90 30 0 30 0 0 2760 0 ;
    END
  END VSS
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2730 270 2690 270 2690 510 2660 510 2660 270 2610 270 2610 510 2580 510 2580 270 2530 270 2530 510 2500 510 2500 270 2450 270 2450 510 2420 510 2420 270 2370 270 2370 510 2340 510 2340 270 2290 270 2290 510 2260 510 2260 270 2210 270 2210 510 2180 510 2180 270 2130 270 2130 510 2100 510 2100 270 2050 270 2050 510 2020 510 2020 270 1970 270 1970 510 1940 510 1940 270 1890 270 1890 510 1860 510 1860 270 1810 270 1810 510 1780 510 1780 270 1730 270 1730 510 1700 510 1700 270 1650 270 1650 510 1620 510 1620 270 1570 270 1570 510 1540 510 1540 270 1490 270 1490 510 1460 510 1460 150 1695 150 1695 130 2495 130 2495 150 2730 150 ;
    END
  END OUT
  PIN IN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.5 612 50.5 702 ;
    END
  END IN1
  PIN IN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20 292 50 382 ;
    END
  END IN2
  OBS
    LAYER M1 ;
      POLYGON 2730 830 2700 830 2700 590 2650 590 2650 830 2620 830 2620 590 2570 590 2570 830 2540 830 2540 590 2490 590 2490 830 2460 830 2460 590 2410 590 2410 830 2380 830 2380 590 2330 590 2330 830 2300 830 2300 590 2250 590 2250 830 2220 830 2220 590 2170 590 2170 830 2140 830 2140 590 2090 590 2090 830 2060 830 2060 590 2010 590 2010 830 1980 830 1980 590 1930 590 1930 830 1900 830 1900 590 1850 590 1850 830 1820 830 1820 590 1770 590 1770 830 1740 830 1740 590 1690 590 1690 830 1660 830 1660 590 1610 590 1610 830 1580 830 1580 590 1530 590 1530 830 1500 830 1500 590 1450 590 1450 830 1420 830 1420 310 1450 310 1450 550 1500 550 1500 310 1530 310 1530 550 1580 550 1580 310 1610 310 1610 550 1660 550 1660 310 1690 310 1690 550 1740 550 1740 310 1770 310 1770 550 1820 550 1820 310 1850 310 1850 550 1900 550 1900 310 1930 310 1930 550 1980 550 1980 310 2010 310 2010 550 2060 550 2060 310 2090 310 2090 550 2140 550 2140 310 2170 310 2170 550 2220 550 2220 310 2250 310 2250 550 2300 550 2300 310 2330 310 2330 550 2380 550 2380 310 2410 310 2410 550 2460 550 2460 310 2490 310 2490 550 2540 550 2540 310 2570 310 2570 550 2620 550 2620 310 2650 310 2650 550 2700 550 2700 310 2730 310 ;
      POLYGON 1380 830 1350 830 1350 590 1300 590 1300 830 1270 830 1270 590 1220 590 1220 830 1190 830 1190 590 1140 590 1140 830 1110 830 1110 590 1060 590 1060 830 1030 830 1030 590 980 590 980 830 950 830 950 590 900 590 900 830 870 830 870 590 820 590 820 830 790 830 790 590 740 590 740 830 710 830 710 590 660 590 660 830 630 830 630 590 580 590 580 830 550 830 550 590 500 590 500 830 470 830 470 590 420 590 420 830 390 830 390 590 340 590 340 830 310 830 310 590 260 590 260 830 230 830 230 590 180 590 180 830 150 830 150 590 100 590 100 830 70 830 70 310 100 310 100 550 150 550 150 310 180 310 180 550 230 550 230 310 260 310 260 550 310 550 310 310 340 310 340 550 390 550 390 310 420 310 420 550 470 550 470 310 500 310 500 550 550 550 550 310 580 310 580 550 630 550 630 310 660 310 660 550 710 550 710 310 740 310 740 550 790 550 790 310 820 310 820 550 870 550 870 310 900 310 900 550 950 550 950 310 980 310 980 550 1030 550 1030 310 1060 310 1060 550 1110 550 1110 310 1140 310 1140 550 1190 550 1190 310 1220 310 1220 550 1270 550 1270 310 1300 310 1300 550 1350 550 1350 310 1380 310 ;
      POLYGON 1340 510 1310 510 1310 270 1260 270 1260 510 1230 510 1230 270 1180 270 1180 510 1150 510 1150 270 1100 270 1100 510 1070 510 1070 270 1020 270 1020 510 990 510 990 270 940 270 940 510 910 510 910 270 860 270 860 510 830 510 830 270 780 270 780 510 750 510 750 270 700 270 700 510 670 510 670 270 620 270 620 510 590 510 590 270 540 270 540 510 510 510 510 270 460 270 460 510 430 510 430 270 380 270 380 510 350 510 350 270 300 270 300 510 270 510 270 270 220 270 220 510 190 510 190 270 140 270 140 510 110 510 110 270 90 270 90 170 890 170 890 190 1340 190 ;
    LAYER Via1 ;
      RECT 1410 240 1420 250 ;
      RECT 1390 240 1400 250 ;
      RECT 1370 240 1380 250 ;
      RECT 1320 240 1330 250 ;
      RECT 1300 240 1310 250 ;
      RECT 1280 240 1290 250 ;
      RECT 950 80 960 90 ;
      RECT 950 130 960 140 ;
      RECT 930 80 940 90 ;
      RECT 930 130 940 140 ;
      RECT 910 80 920 90 ;
      RECT 910 130 920 140 ;
      RECT 30.5 622 40.5 632 ;
      RECT 30.5 642 40.5 652 ;
      RECT 30.5 662 40.5 672 ;
      RECT 30.5 682 40.5 692 ;
      RECT 30 302 40 312 ;
      RECT 30 322 40 332 ;
      RECT 30 342 40 352 ;
      RECT 30 362 40 372 ;
    LAYER M2 ;
      RECT 1270 230 1430 260 ;
  END
END NOR2D8

END LIBRARY
