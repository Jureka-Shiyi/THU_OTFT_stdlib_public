* SPICE NETLIST
***************************************

.SUBCKT BOUNDARY_LEFT
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
